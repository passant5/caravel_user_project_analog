magic
tech sky130A
magscale 1 2
timestamp 1684745564
<< obsli1 >>
rect 1104 2159 582820 701777
<< obsm1 >>
rect 566 1368 582990 702296
<< metal2 >>
rect 1278 703520 1390 704960
rect 5142 703520 5254 704960
rect 9006 703520 9118 704960
rect 12870 703520 12982 704960
rect 16090 703520 16202 704960
rect 19954 703520 20066 704960
rect 23818 703520 23930 704960
rect 27682 703520 27794 704960
rect 31546 703520 31658 704960
rect 35410 703520 35522 704960
rect 39274 703520 39386 704960
rect 43138 703520 43250 704960
rect 47002 703520 47114 704960
rect 50866 703520 50978 704960
rect 54730 703520 54842 704960
rect 58594 703520 58706 704960
rect 62458 703520 62570 704960
rect 66322 703520 66434 704960
rect 70186 703520 70298 704960
rect 73406 703520 73518 704960
rect 77270 703520 77382 704960
rect 81134 703520 81246 704960
rect 84998 703520 85110 704960
rect 88862 703520 88974 704960
rect 92726 703520 92838 704960
rect 96590 703520 96702 704960
rect 100454 703520 100566 704960
rect 104318 703520 104430 704960
rect 108182 703520 108294 704960
rect 112046 703520 112158 704960
rect 115910 703520 116022 704960
rect 119774 703520 119886 704960
rect 123638 703520 123750 704960
rect 127502 703520 127614 704960
rect 130722 703520 130834 704960
rect 134586 703520 134698 704960
rect 138450 703520 138562 704960
rect 142314 703520 142426 704960
rect 146178 703520 146290 704960
rect 150042 703520 150154 704960
rect 153906 703520 154018 704960
rect 157770 703520 157882 704960
rect 161634 703520 161746 704960
rect 165498 703520 165610 704960
rect 169362 703520 169474 704960
rect 173226 703520 173338 704960
rect 177090 703520 177202 704960
rect 180954 703520 181066 704960
rect 184818 703520 184930 704960
rect 188038 703520 188150 704960
rect 191902 703520 192014 704960
rect 195766 703520 195878 704960
rect 199630 703520 199742 704960
rect 203494 703520 203606 704960
rect 207358 703520 207470 704960
rect 211222 703520 211334 704960
rect 215086 703520 215198 704960
rect 218950 703520 219062 704960
rect 222814 703520 222926 704960
rect 226678 703520 226790 704960
rect 230542 703520 230654 704960
rect 234406 703520 234518 704960
rect 238270 703520 238382 704960
rect 242134 703520 242246 704960
rect 245354 703520 245466 704960
rect 249218 703520 249330 704960
rect 253082 703520 253194 704960
rect 256946 703520 257058 704960
rect 260810 703520 260922 704960
rect 264674 703520 264786 704960
rect 268538 703520 268650 704960
rect 272402 703520 272514 704960
rect 276266 703520 276378 704960
rect 280130 703520 280242 704960
rect 283994 703520 284106 704960
rect 287858 703520 287970 704960
rect 291722 703520 291834 704960
rect 295586 703520 295698 704960
rect 299450 703520 299562 704960
rect 302670 703520 302782 704960
rect 306534 703520 306646 704960
rect 310398 703520 310510 704960
rect 314262 703520 314374 704960
rect 318126 703520 318238 704960
rect 321990 703520 322102 704960
rect 325854 703520 325966 704960
rect 329718 703520 329830 704960
rect 333582 703520 333694 704960
rect 337446 703520 337558 704960
rect 341310 703520 341422 704960
rect 345174 703520 345286 704960
rect 349038 703520 349150 704960
rect 352902 703520 353014 704960
rect 356122 703520 356234 704960
rect 359986 703520 360098 704960
rect 363850 703520 363962 704960
rect 367714 703520 367826 704960
rect 371578 703520 371690 704960
rect 375442 703520 375554 704960
rect 379306 703520 379418 704960
rect 383170 703520 383282 704960
rect 387034 703520 387146 704960
rect 390898 703520 391010 704960
rect 394762 703520 394874 704960
rect 398626 703520 398738 704960
rect 402490 703520 402602 704960
rect 406354 703520 406466 704960
rect 410218 703520 410330 704960
rect 413438 703520 413550 704960
rect 417302 703520 417414 704960
rect 421166 703520 421278 704960
rect 425030 703520 425142 704960
rect 428894 703520 429006 704960
rect 432758 703520 432870 704960
rect 436622 703520 436734 704960
rect 440486 703520 440598 704960
rect 444350 703520 444462 704960
rect 448214 703520 448326 704960
rect 452078 703520 452190 704960
rect 455942 703520 456054 704960
rect 459806 703520 459918 704960
rect 463670 703520 463782 704960
rect 467534 703520 467646 704960
rect 470754 703520 470866 704960
rect 474618 703520 474730 704960
rect 478482 703520 478594 704960
rect 482346 703520 482458 704960
rect 486210 703520 486322 704960
rect 490074 703520 490186 704960
rect 493938 703520 494050 704960
rect 497802 703520 497914 704960
rect 501666 703520 501778 704960
rect 505530 703520 505642 704960
rect 509394 703520 509506 704960
rect 513258 703520 513370 704960
rect 517122 703520 517234 704960
rect 520986 703520 521098 704960
rect 524850 703520 524962 704960
rect 528070 703520 528182 704960
rect 531934 703520 532046 704960
rect 535798 703520 535910 704960
rect 539662 703520 539774 704960
rect 543526 703520 543638 704960
rect 547390 703520 547502 704960
rect 551254 703520 551366 704960
rect 555118 703520 555230 704960
rect 558982 703520 559094 704960
rect 562846 703520 562958 704960
rect 566710 703520 566822 704960
rect 570574 703520 570686 704960
rect 574438 703520 574550 704960
rect 578302 703520 578414 704960
rect 582166 703520 582278 704960
rect -10 -960 102 480
rect 3210 -960 3322 480
rect 7074 -960 7186 480
rect 10938 -960 11050 480
rect 14802 -960 14914 480
rect 18666 -960 18778 480
rect 22530 -960 22642 480
rect 26394 -960 26506 480
rect 30258 -960 30370 480
rect 34122 -960 34234 480
rect 37986 -960 38098 480
rect 41850 -960 41962 480
rect 45714 -960 45826 480
rect 49578 -960 49690 480
rect 53442 -960 53554 480
rect 56662 -960 56774 480
rect 60526 -960 60638 480
rect 64390 -960 64502 480
rect 68254 -960 68366 480
rect 72118 -960 72230 480
rect 75982 -960 76094 480
rect 79846 -960 79958 480
rect 83710 -960 83822 480
rect 87574 -960 87686 480
rect 91438 -960 91550 480
rect 95302 -960 95414 480
rect 99166 -960 99278 480
rect 103030 -960 103142 480
rect 106894 -960 107006 480
rect 110758 -960 110870 480
rect 113978 -960 114090 480
rect 117842 -960 117954 480
rect 121706 -960 121818 480
rect 125570 -960 125682 480
rect 129434 -960 129546 480
rect 133298 -960 133410 480
rect 137162 -960 137274 480
rect 141026 -960 141138 480
rect 144890 -960 145002 480
rect 148754 -960 148866 480
rect 152618 -960 152730 480
rect 156482 -960 156594 480
rect 160346 -960 160458 480
rect 164210 -960 164322 480
rect 168074 -960 168186 480
rect 171294 -960 171406 480
rect 175158 -960 175270 480
rect 179022 -960 179134 480
rect 182886 -960 182998 480
rect 186750 -960 186862 480
rect 190614 -960 190726 480
rect 194478 -960 194590 480
rect 198342 -960 198454 480
rect 202206 -960 202318 480
rect 206070 -960 206182 480
rect 209934 -960 210046 480
rect 213798 -960 213910 480
rect 217662 -960 217774 480
rect 221526 -960 221638 480
rect 225390 -960 225502 480
rect 228610 -960 228722 480
rect 232474 -960 232586 480
rect 236338 -960 236450 480
rect 240202 -960 240314 480
rect 244066 -960 244178 480
rect 247930 -960 248042 480
rect 251794 -960 251906 480
rect 255658 -960 255770 480
rect 259522 -960 259634 480
rect 263386 -960 263498 480
rect 267250 -960 267362 480
rect 271114 -960 271226 480
rect 274978 -960 275090 480
rect 278842 -960 278954 480
rect 282706 -960 282818 480
rect 285926 -960 286038 480
rect 289790 -960 289902 480
rect 293654 -960 293766 480
rect 297518 -960 297630 480
rect 301382 -960 301494 480
rect 305246 -960 305358 480
rect 309110 -960 309222 480
rect 312974 -960 313086 480
rect 316838 -960 316950 480
rect 320702 -960 320814 480
rect 324566 -960 324678 480
rect 328430 -960 328542 480
rect 332294 -960 332406 480
rect 336158 -960 336270 480
rect 340022 -960 340134 480
rect 343242 -960 343354 480
rect 347106 -960 347218 480
rect 350970 -960 351082 480
rect 354834 -960 354946 480
rect 358698 -960 358810 480
rect 362562 -960 362674 480
rect 366426 -960 366538 480
rect 370290 -960 370402 480
rect 374154 -960 374266 480
rect 378018 -960 378130 480
rect 381882 -960 381994 480
rect 385746 -960 385858 480
rect 389610 -960 389722 480
rect 393474 -960 393586 480
rect 397338 -960 397450 480
rect 400558 -960 400670 480
rect 404422 -960 404534 480
rect 408286 -960 408398 480
rect 412150 -960 412262 480
rect 416014 -960 416126 480
rect 419878 -960 419990 480
rect 423742 -960 423854 480
rect 427606 -960 427718 480
rect 431470 -960 431582 480
rect 435334 -960 435446 480
rect 439198 -960 439310 480
rect 443062 -960 443174 480
rect 446926 -960 447038 480
rect 450790 -960 450902 480
rect 454654 -960 454766 480
rect 457874 -960 457986 480
rect 461738 -960 461850 480
rect 465602 -960 465714 480
rect 469466 -960 469578 480
rect 473330 -960 473442 480
rect 477194 -960 477306 480
rect 481058 -960 481170 480
rect 484922 -960 485034 480
rect 488786 -960 488898 480
rect 492650 -960 492762 480
rect 496514 -960 496626 480
rect 500378 -960 500490 480
rect 504242 -960 504354 480
rect 508106 -960 508218 480
rect 511326 -960 511438 480
rect 515190 -960 515302 480
rect 519054 -960 519166 480
rect 522918 -960 523030 480
rect 526782 -960 526894 480
rect 530646 -960 530758 480
rect 534510 -960 534622 480
rect 538374 -960 538486 480
rect 542238 -960 542350 480
rect 546102 -960 546214 480
rect 549966 -960 550078 480
rect 553830 -960 553942 480
rect 557694 -960 557806 480
rect 561558 -960 561670 480
rect 565422 -960 565534 480
rect 568642 -960 568754 480
rect 572506 -960 572618 480
rect 576370 -960 576482 480
rect 580234 -960 580346 480
<< obsm2 >>
rect 18 703464 1222 703610
rect 1446 703464 5086 703610
rect 5310 703464 8950 703610
rect 9174 703464 12814 703610
rect 13038 703464 16034 703610
rect 16258 703464 19898 703610
rect 20122 703464 23762 703610
rect 23986 703464 27626 703610
rect 27850 703464 31490 703610
rect 31714 703464 35354 703610
rect 35578 703464 39218 703610
rect 39442 703464 43082 703610
rect 43306 703464 46946 703610
rect 47170 703464 50810 703610
rect 51034 703464 54674 703610
rect 54898 703464 58538 703610
rect 58762 703464 62402 703610
rect 62626 703464 66266 703610
rect 66490 703464 70130 703610
rect 70354 703464 73350 703610
rect 73574 703464 77214 703610
rect 77438 703464 81078 703610
rect 81302 703464 84942 703610
rect 85166 703464 88806 703610
rect 89030 703464 92670 703610
rect 92894 703464 96534 703610
rect 96758 703464 100398 703610
rect 100622 703464 104262 703610
rect 104486 703464 108126 703610
rect 108350 703464 111990 703610
rect 112214 703464 115854 703610
rect 116078 703464 119718 703610
rect 119942 703464 123582 703610
rect 123806 703464 127446 703610
rect 127670 703464 130666 703610
rect 130890 703464 134530 703610
rect 134754 703464 138394 703610
rect 138618 703464 142258 703610
rect 142482 703464 146122 703610
rect 146346 703464 149986 703610
rect 150210 703464 153850 703610
rect 154074 703464 157714 703610
rect 157938 703464 161578 703610
rect 161802 703464 165442 703610
rect 165666 703464 169306 703610
rect 169530 703464 173170 703610
rect 173394 703464 177034 703610
rect 177258 703464 180898 703610
rect 181122 703464 184762 703610
rect 184986 703464 187982 703610
rect 188206 703464 191846 703610
rect 192070 703464 195710 703610
rect 195934 703464 199574 703610
rect 199798 703464 203438 703610
rect 203662 703464 207302 703610
rect 207526 703464 211166 703610
rect 211390 703464 215030 703610
rect 215254 703464 218894 703610
rect 219118 703464 222758 703610
rect 222982 703464 226622 703610
rect 226846 703464 230486 703610
rect 230710 703464 234350 703610
rect 234574 703464 238214 703610
rect 238438 703464 242078 703610
rect 242302 703464 245298 703610
rect 245522 703464 249162 703610
rect 249386 703464 253026 703610
rect 253250 703464 256890 703610
rect 257114 703464 260754 703610
rect 260978 703464 264618 703610
rect 264842 703464 268482 703610
rect 268706 703464 272346 703610
rect 272570 703464 276210 703610
rect 276434 703464 280074 703610
rect 280298 703464 283938 703610
rect 284162 703464 287802 703610
rect 288026 703464 291666 703610
rect 291890 703464 295530 703610
rect 295754 703464 299394 703610
rect 299618 703464 302614 703610
rect 302838 703464 306478 703610
rect 306702 703464 310342 703610
rect 310566 703464 314206 703610
rect 314430 703464 318070 703610
rect 318294 703464 321934 703610
rect 322158 703464 325798 703610
rect 326022 703464 329662 703610
rect 329886 703464 333526 703610
rect 333750 703464 337390 703610
rect 337614 703464 341254 703610
rect 341478 703464 345118 703610
rect 345342 703464 348982 703610
rect 349206 703464 352846 703610
rect 353070 703464 356066 703610
rect 356290 703464 359930 703610
rect 360154 703464 363794 703610
rect 364018 703464 367658 703610
rect 367882 703464 371522 703610
rect 371746 703464 375386 703610
rect 375610 703464 379250 703610
rect 379474 703464 383114 703610
rect 383338 703464 386978 703610
rect 387202 703464 390842 703610
rect 391066 703464 394706 703610
rect 394930 703464 398570 703610
rect 398794 703464 402434 703610
rect 402658 703464 406298 703610
rect 406522 703464 410162 703610
rect 410386 703464 413382 703610
rect 413606 703464 417246 703610
rect 417470 703464 421110 703610
rect 421334 703464 424974 703610
rect 425198 703464 428838 703610
rect 429062 703464 432702 703610
rect 432926 703464 436566 703610
rect 436790 703464 440430 703610
rect 440654 703464 444294 703610
rect 444518 703464 448158 703610
rect 448382 703464 452022 703610
rect 452246 703464 455886 703610
rect 456110 703464 459750 703610
rect 459974 703464 463614 703610
rect 463838 703464 467478 703610
rect 467702 703464 470698 703610
rect 470922 703464 474562 703610
rect 474786 703464 478426 703610
rect 478650 703464 482290 703610
rect 482514 703464 486154 703610
rect 486378 703464 490018 703610
rect 490242 703464 493882 703610
rect 494106 703464 497746 703610
rect 497970 703464 501610 703610
rect 501834 703464 505474 703610
rect 505698 703464 509338 703610
rect 509562 703464 513202 703610
rect 513426 703464 517066 703610
rect 517290 703464 520930 703610
rect 521154 703464 524794 703610
rect 525018 703464 528014 703610
rect 528238 703464 531878 703610
rect 532102 703464 535742 703610
rect 535966 703464 539606 703610
rect 539830 703464 543470 703610
rect 543694 703464 547334 703610
rect 547558 703464 551198 703610
rect 551422 703464 555062 703610
rect 555286 703464 558926 703610
rect 559150 703464 562790 703610
rect 563014 703464 566654 703610
rect 566878 703464 570518 703610
rect 570742 703464 574382 703610
rect 574606 703464 578246 703610
rect 578470 703464 582110 703610
rect 582334 703464 582984 703610
rect 18 536 582984 703464
rect 158 31 3154 536
rect 3378 31 7018 536
rect 7242 31 10882 536
rect 11106 31 14746 536
rect 14970 31 18610 536
rect 18834 31 22474 536
rect 22698 31 26338 536
rect 26562 31 30202 536
rect 30426 31 34066 536
rect 34290 31 37930 536
rect 38154 31 41794 536
rect 42018 31 45658 536
rect 45882 31 49522 536
rect 49746 31 53386 536
rect 53610 31 56606 536
rect 56830 31 60470 536
rect 60694 31 64334 536
rect 64558 31 68198 536
rect 68422 31 72062 536
rect 72286 31 75926 536
rect 76150 31 79790 536
rect 80014 31 83654 536
rect 83878 31 87518 536
rect 87742 31 91382 536
rect 91606 31 95246 536
rect 95470 31 99110 536
rect 99334 31 102974 536
rect 103198 31 106838 536
rect 107062 31 110702 536
rect 110926 31 113922 536
rect 114146 31 117786 536
rect 118010 31 121650 536
rect 121874 31 125514 536
rect 125738 31 129378 536
rect 129602 31 133242 536
rect 133466 31 137106 536
rect 137330 31 140970 536
rect 141194 31 144834 536
rect 145058 31 148698 536
rect 148922 31 152562 536
rect 152786 31 156426 536
rect 156650 31 160290 536
rect 160514 31 164154 536
rect 164378 31 168018 536
rect 168242 31 171238 536
rect 171462 31 175102 536
rect 175326 31 178966 536
rect 179190 31 182830 536
rect 183054 31 186694 536
rect 186918 31 190558 536
rect 190782 31 194422 536
rect 194646 31 198286 536
rect 198510 31 202150 536
rect 202374 31 206014 536
rect 206238 31 209878 536
rect 210102 31 213742 536
rect 213966 31 217606 536
rect 217830 31 221470 536
rect 221694 31 225334 536
rect 225558 31 228554 536
rect 228778 31 232418 536
rect 232642 31 236282 536
rect 236506 31 240146 536
rect 240370 31 244010 536
rect 244234 31 247874 536
rect 248098 31 251738 536
rect 251962 31 255602 536
rect 255826 31 259466 536
rect 259690 31 263330 536
rect 263554 31 267194 536
rect 267418 31 271058 536
rect 271282 31 274922 536
rect 275146 31 278786 536
rect 279010 31 282650 536
rect 282874 31 285870 536
rect 286094 31 289734 536
rect 289958 31 293598 536
rect 293822 31 297462 536
rect 297686 31 301326 536
rect 301550 31 305190 536
rect 305414 31 309054 536
rect 309278 31 312918 536
rect 313142 31 316782 536
rect 317006 31 320646 536
rect 320870 31 324510 536
rect 324734 31 328374 536
rect 328598 31 332238 536
rect 332462 31 336102 536
rect 336326 31 339966 536
rect 340190 31 343186 536
rect 343410 31 347050 536
rect 347274 31 350914 536
rect 351138 31 354778 536
rect 355002 31 358642 536
rect 358866 31 362506 536
rect 362730 31 366370 536
rect 366594 31 370234 536
rect 370458 31 374098 536
rect 374322 31 377962 536
rect 378186 31 381826 536
rect 382050 31 385690 536
rect 385914 31 389554 536
rect 389778 31 393418 536
rect 393642 31 397282 536
rect 397506 31 400502 536
rect 400726 31 404366 536
rect 404590 31 408230 536
rect 408454 31 412094 536
rect 412318 31 415958 536
rect 416182 31 419822 536
rect 420046 31 423686 536
rect 423910 31 427550 536
rect 427774 31 431414 536
rect 431638 31 435278 536
rect 435502 31 439142 536
rect 439366 31 443006 536
rect 443230 31 446870 536
rect 447094 31 450734 536
rect 450958 31 454598 536
rect 454822 31 457818 536
rect 458042 31 461682 536
rect 461906 31 465546 536
rect 465770 31 469410 536
rect 469634 31 473274 536
rect 473498 31 477138 536
rect 477362 31 481002 536
rect 481226 31 484866 536
rect 485090 31 488730 536
rect 488954 31 492594 536
rect 492818 31 496458 536
rect 496682 31 500322 536
rect 500546 31 504186 536
rect 504410 31 508050 536
rect 508274 31 511270 536
rect 511494 31 515134 536
rect 515358 31 518998 536
rect 519222 31 522862 536
rect 523086 31 526726 536
rect 526950 31 530590 536
rect 530814 31 534454 536
rect 534678 31 538318 536
rect 538542 31 542182 536
rect 542406 31 546046 536
rect 546270 31 549910 536
rect 550134 31 553774 536
rect 553998 31 557638 536
rect 557862 31 561502 536
rect 561726 31 565366 536
rect 565590 31 568586 536
rect 568810 31 572450 536
rect 572674 31 576314 536
rect 576538 31 580178 536
rect 580402 31 582984 536
<< metal3 >>
rect 583520 702388 584960 702628
rect -960 701708 480 701948
rect 583520 698308 584960 698548
rect -960 697628 480 697868
rect 583520 694228 584960 694468
rect -960 693548 480 693788
rect 583520 690148 584960 690388
rect -960 689468 480 689708
rect 583520 686068 584960 686308
rect -960 685388 480 685628
rect 583520 681988 584960 682228
rect -960 681308 480 681548
rect 583520 677908 584960 678148
rect -960 677228 480 677468
rect 583520 673828 584960 674068
rect -960 673148 480 673388
rect 583520 669748 584960 669988
rect -960 669068 480 669308
rect 583520 665668 584960 665908
rect -960 664988 480 665228
rect 583520 661588 584960 661828
rect -960 660908 480 661148
rect -960 657508 480 657748
rect 583520 657508 584960 657748
rect -960 653428 480 653668
rect 583520 653428 584960 653668
rect -960 649348 480 649588
rect 583520 649348 584960 649588
rect -960 645268 480 645508
rect 583520 645268 584960 645508
rect 583520 641868 584960 642108
rect -960 641188 480 641428
rect 583520 637788 584960 638028
rect -960 637108 480 637348
rect 583520 633708 584960 633948
rect -960 633028 480 633268
rect 583520 629628 584960 629868
rect -960 628948 480 629188
rect 583520 625548 584960 625788
rect -960 624868 480 625108
rect 583520 621468 584960 621708
rect -960 620788 480 621028
rect 583520 617388 584960 617628
rect -960 616708 480 616948
rect 583520 613308 584960 613548
rect -960 612628 480 612868
rect 583520 609228 584960 609468
rect -960 608548 480 608788
rect 583520 605148 584960 605388
rect -960 604468 480 604708
rect 583520 601068 584960 601308
rect -960 600388 480 600628
rect -960 596988 480 597228
rect 583520 596988 584960 597228
rect -960 592908 480 593148
rect 583520 592908 584960 593148
rect -960 588828 480 589068
rect 583520 588828 584960 589068
rect -960 584748 480 584988
rect 583520 584748 584960 584988
rect 583520 581348 584960 581588
rect -960 580668 480 580908
rect 583520 577268 584960 577508
rect -960 576588 480 576828
rect 583520 573188 584960 573428
rect -960 572508 480 572748
rect 583520 569108 584960 569348
rect -960 568428 480 568668
rect 583520 565028 584960 565268
rect -960 564348 480 564588
rect 583520 560948 584960 561188
rect -960 560268 480 560508
rect 583520 556868 584960 557108
rect -960 556188 480 556428
rect 583520 552788 584960 553028
rect -960 552108 480 552348
rect 583520 548708 584960 548948
rect -960 548028 480 548268
rect 583520 544628 584960 544868
rect -960 543948 480 544188
rect 583520 540548 584960 540788
rect -960 539868 480 540108
rect -960 536468 480 536708
rect 583520 536468 584960 536708
rect -960 532388 480 532628
rect 583520 532388 584960 532628
rect -960 528308 480 528548
rect 583520 528308 584960 528548
rect -960 524228 480 524468
rect 583520 524228 584960 524468
rect 583520 520828 584960 521068
rect -960 520148 480 520388
rect 583520 516748 584960 516988
rect -960 516068 480 516308
rect 583520 512668 584960 512908
rect -960 511988 480 512228
rect 583520 508588 584960 508828
rect -960 507908 480 508148
rect 583520 504508 584960 504748
rect -960 503828 480 504068
rect 583520 500428 584960 500668
rect -960 499748 480 499988
rect 583520 496348 584960 496588
rect -960 495668 480 495908
rect 583520 492268 584960 492508
rect -960 491588 480 491828
rect 583520 488188 584960 488428
rect -960 487508 480 487748
rect 583520 484108 584960 484348
rect -960 483428 480 483668
rect -960 480028 480 480268
rect 583520 480028 584960 480268
rect -960 475948 480 476188
rect 583520 475948 584960 476188
rect -960 471868 480 472108
rect 583520 471868 584960 472108
rect -960 467788 480 468028
rect 583520 467788 584960 468028
rect -960 463708 480 463948
rect 583520 463708 584960 463948
rect 583520 460308 584960 460548
rect -960 459628 480 459868
rect 583520 456228 584960 456468
rect -960 455548 480 455788
rect 583520 452148 584960 452388
rect -960 451468 480 451708
rect 583520 448068 584960 448308
rect -960 447388 480 447628
rect 583520 443988 584960 444228
rect -960 443308 480 443548
rect 583520 439908 584960 440148
rect -960 439228 480 439468
rect 583520 435828 584960 436068
rect -960 435148 480 435388
rect 583520 431748 584960 431988
rect -960 431068 480 431308
rect 583520 427668 584960 427908
rect -960 426988 480 427228
rect 583520 423588 584960 423828
rect -960 422908 480 423148
rect -960 419508 480 419748
rect 583520 419508 584960 419748
rect -960 415428 480 415668
rect 583520 415428 584960 415668
rect -960 411348 480 411588
rect 583520 411348 584960 411588
rect -960 407268 480 407508
rect 583520 407268 584960 407508
rect 583520 403868 584960 404108
rect -960 403188 480 403428
rect 583520 399788 584960 400028
rect -960 399108 480 399348
rect 583520 395708 584960 395948
rect -960 395028 480 395268
rect 583520 391628 584960 391868
rect -960 390948 480 391188
rect 583520 387548 584960 387788
rect -960 386868 480 387108
rect 583520 383468 584960 383708
rect -960 382788 480 383028
rect 583520 379388 584960 379628
rect -960 378708 480 378948
rect 583520 375308 584960 375548
rect -960 374628 480 374868
rect 583520 371228 584960 371468
rect -960 370548 480 370788
rect 583520 367148 584960 367388
rect -960 366468 480 366708
rect 583520 363068 584960 363308
rect -960 362388 480 362628
rect -960 358988 480 359228
rect 583520 358988 584960 359228
rect -960 354908 480 355148
rect 583520 354908 584960 355148
rect -960 350828 480 351068
rect 583520 350828 584960 351068
rect -960 346748 480 346988
rect 583520 346748 584960 346988
rect 583520 343348 584960 343588
rect -960 342668 480 342908
rect 583520 339268 584960 339508
rect -960 338588 480 338828
rect 583520 335188 584960 335428
rect -960 334508 480 334748
rect 583520 331108 584960 331348
rect -960 330428 480 330668
rect 583520 327028 584960 327268
rect -960 326348 480 326588
rect 583520 322948 584960 323188
rect -960 322268 480 322508
rect 583520 318868 584960 319108
rect -960 318188 480 318428
rect 583520 314788 584960 315028
rect -960 314108 480 314348
rect 583520 310708 584960 310948
rect -960 310028 480 310268
rect 583520 306628 584960 306868
rect -960 305948 480 306188
rect 583520 302548 584960 302788
rect -960 301868 480 302108
rect -960 298468 480 298708
rect 583520 298468 584960 298708
rect -960 294388 480 294628
rect 583520 294388 584960 294628
rect -960 290308 480 290548
rect 583520 290308 584960 290548
rect -960 286228 480 286468
rect 583520 286228 584960 286468
rect 583520 282828 584960 283068
rect -960 282148 480 282388
rect 583520 278748 584960 278988
rect -960 278068 480 278308
rect 583520 274668 584960 274908
rect -960 273988 480 274228
rect 583520 270588 584960 270828
rect -960 269908 480 270148
rect 583520 266508 584960 266748
rect -960 265828 480 266068
rect 583520 262428 584960 262668
rect -960 261748 480 261988
rect 583520 258348 584960 258588
rect -960 257668 480 257908
rect 583520 254268 584960 254508
rect -960 253588 480 253828
rect 583520 250188 584960 250428
rect -960 249508 480 249748
rect 583520 246108 584960 246348
rect -960 245428 480 245668
rect 583520 242028 584960 242268
rect -960 241348 480 241588
rect -960 237948 480 238188
rect 583520 237948 584960 238188
rect -960 233868 480 234108
rect 583520 233868 584960 234108
rect -960 229788 480 230028
rect 583520 229788 584960 230028
rect -960 225708 480 225948
rect 583520 225708 584960 225948
rect 583520 222308 584960 222548
rect -960 221628 480 221868
rect 583520 218228 584960 218468
rect -960 217548 480 217788
rect 583520 214148 584960 214388
rect -960 213468 480 213708
rect 583520 210068 584960 210308
rect -960 209388 480 209628
rect 583520 205988 584960 206228
rect -960 205308 480 205548
rect 583520 201908 584960 202148
rect -960 201228 480 201468
rect 583520 197828 584960 198068
rect -960 197148 480 197388
rect 583520 193748 584960 193988
rect -960 193068 480 193308
rect 583520 189668 584960 189908
rect -960 188988 480 189228
rect 583520 185588 584960 185828
rect -960 184908 480 185148
rect 583520 181508 584960 181748
rect -960 180828 480 181068
rect -960 177428 480 177668
rect 583520 177428 584960 177668
rect -960 173348 480 173588
rect 583520 173348 584960 173588
rect -960 169268 480 169508
rect 583520 169268 584960 169508
rect -960 165188 480 165428
rect 583520 165188 584960 165428
rect 583520 161788 584960 162028
rect -960 161108 480 161348
rect 583520 157708 584960 157948
rect -960 157028 480 157268
rect 583520 153628 584960 153868
rect -960 152948 480 153188
rect 583520 149548 584960 149788
rect -960 148868 480 149108
rect 583520 145468 584960 145708
rect -960 144788 480 145028
rect 583520 141388 584960 141628
rect -960 140708 480 140948
rect 583520 137308 584960 137548
rect -960 136628 480 136868
rect 583520 133228 584960 133468
rect -960 132548 480 132788
rect 583520 129148 584960 129388
rect -960 128468 480 128708
rect 583520 125068 584960 125308
rect -960 124388 480 124628
rect 583520 120988 584960 121228
rect -960 120308 480 120548
rect -960 116908 480 117148
rect 583520 116908 584960 117148
rect -960 112828 480 113068
rect 583520 112828 584960 113068
rect -960 108748 480 108988
rect 583520 108748 584960 108988
rect -960 104668 480 104908
rect 583520 104668 584960 104908
rect 583520 101268 584960 101508
rect -960 100588 480 100828
rect 583520 97188 584960 97428
rect -960 96508 480 96748
rect 583520 93108 584960 93348
rect -960 92428 480 92668
rect 583520 89028 584960 89268
rect -960 88348 480 88588
rect 583520 84948 584960 85188
rect -960 84268 480 84508
rect 583520 80868 584960 81108
rect -960 80188 480 80428
rect 583520 76788 584960 77028
rect -960 76108 480 76348
rect 583520 72708 584960 72948
rect -960 72028 480 72268
rect 583520 68628 584960 68868
rect -960 67948 480 68188
rect 583520 64548 584960 64788
rect -960 63868 480 64108
rect 583520 60468 584960 60708
rect -960 59788 480 60028
rect -960 56388 480 56628
rect 583520 56388 584960 56628
rect -960 52308 480 52548
rect 583520 52308 584960 52548
rect -960 48228 480 48468
rect 583520 48228 584960 48468
rect -960 44148 480 44388
rect 583520 44148 584960 44388
rect 583520 40748 584960 40988
rect -960 40068 480 40308
rect 583520 36668 584960 36908
rect -960 35988 480 36228
rect 583520 32588 584960 32828
rect -960 31908 480 32148
rect 583520 28508 584960 28748
rect -960 27828 480 28068
rect 583520 24428 584960 24668
rect -960 23748 480 23988
rect 583520 20348 584960 20588
rect -960 19668 480 19908
rect 583520 16268 584960 16508
rect -960 15588 480 15828
rect 583520 12188 584960 12428
rect -960 11508 480 11748
rect 583520 8108 584960 8348
rect -960 7428 480 7668
rect 583520 4028 584960 4268
rect -960 3348 480 3588
rect 583520 -52 584960 188
<< obsm3 >>
rect 13 702308 583440 702541
rect 13 702028 583586 702308
rect 560 701628 583586 702028
rect 13 698628 583586 701628
rect 13 698228 583440 698628
rect 13 697948 583586 698228
rect 560 697548 583586 697948
rect 13 694548 583586 697548
rect 13 694148 583440 694548
rect 13 693868 583586 694148
rect 560 693468 583586 693868
rect 13 690468 583586 693468
rect 13 690068 583440 690468
rect 13 689788 583586 690068
rect 560 689388 583586 689788
rect 13 686388 583586 689388
rect 13 685988 583440 686388
rect 13 685708 583586 685988
rect 560 685308 583586 685708
rect 13 682308 583586 685308
rect 13 681908 583440 682308
rect 13 681628 583586 681908
rect 560 681228 583586 681628
rect 13 678228 583586 681228
rect 13 677828 583440 678228
rect 13 677548 583586 677828
rect 560 677148 583586 677548
rect 13 674148 583586 677148
rect 13 673748 583440 674148
rect 13 673468 583586 673748
rect 560 673068 583586 673468
rect 13 670068 583586 673068
rect 13 669668 583440 670068
rect 13 669388 583586 669668
rect 560 668988 583586 669388
rect 13 665988 583586 668988
rect 13 665588 583440 665988
rect 13 665308 583586 665588
rect 560 664908 583586 665308
rect 13 661908 583586 664908
rect 13 661508 583440 661908
rect 13 661228 583586 661508
rect 560 660828 583586 661228
rect 13 657828 583586 660828
rect 560 657428 583440 657828
rect 13 653748 583586 657428
rect 560 653348 583440 653748
rect 13 649668 583586 653348
rect 560 649268 583440 649668
rect 13 645588 583586 649268
rect 560 645188 583440 645588
rect 13 642188 583586 645188
rect 13 641788 583440 642188
rect 13 641508 583586 641788
rect 560 641108 583586 641508
rect 13 638108 583586 641108
rect 13 637708 583440 638108
rect 13 637428 583586 637708
rect 560 637028 583586 637428
rect 13 634028 583586 637028
rect 13 633628 583440 634028
rect 13 633348 583586 633628
rect 560 632948 583586 633348
rect 13 629948 583586 632948
rect 13 629548 583440 629948
rect 13 629268 583586 629548
rect 560 628868 583586 629268
rect 13 625868 583586 628868
rect 13 625468 583440 625868
rect 13 625188 583586 625468
rect 560 624788 583586 625188
rect 13 621788 583586 624788
rect 13 621388 583440 621788
rect 13 621108 583586 621388
rect 560 620708 583586 621108
rect 13 617708 583586 620708
rect 13 617308 583440 617708
rect 13 617028 583586 617308
rect 560 616628 583586 617028
rect 13 613628 583586 616628
rect 13 613228 583440 613628
rect 13 612948 583586 613228
rect 560 612548 583586 612948
rect 13 609548 583586 612548
rect 13 609148 583440 609548
rect 13 608868 583586 609148
rect 560 608468 583586 608868
rect 13 605468 583586 608468
rect 13 605068 583440 605468
rect 13 604788 583586 605068
rect 560 604388 583586 604788
rect 13 601388 583586 604388
rect 13 600988 583440 601388
rect 13 600708 583586 600988
rect 560 600308 583586 600708
rect 13 597308 583586 600308
rect 560 596908 583440 597308
rect 13 593228 583586 596908
rect 560 592828 583440 593228
rect 13 589148 583586 592828
rect 560 588748 583440 589148
rect 13 585068 583586 588748
rect 560 584668 583440 585068
rect 13 581668 583586 584668
rect 13 581268 583440 581668
rect 13 580988 583586 581268
rect 560 580588 583586 580988
rect 13 577588 583586 580588
rect 13 577188 583440 577588
rect 13 576908 583586 577188
rect 560 576508 583586 576908
rect 13 573508 583586 576508
rect 13 573108 583440 573508
rect 13 572828 583586 573108
rect 560 572428 583586 572828
rect 13 569428 583586 572428
rect 13 569028 583440 569428
rect 13 568748 583586 569028
rect 560 568348 583586 568748
rect 13 565348 583586 568348
rect 13 564948 583440 565348
rect 13 564668 583586 564948
rect 560 564268 583586 564668
rect 13 561268 583586 564268
rect 13 560868 583440 561268
rect 13 560588 583586 560868
rect 560 560188 583586 560588
rect 13 557188 583586 560188
rect 13 556788 583440 557188
rect 13 556508 583586 556788
rect 560 556108 583586 556508
rect 13 553108 583586 556108
rect 13 552708 583440 553108
rect 13 552428 583586 552708
rect 560 552028 583586 552428
rect 13 549028 583586 552028
rect 13 548628 583440 549028
rect 13 548348 583586 548628
rect 560 547948 583586 548348
rect 13 544948 583586 547948
rect 13 544548 583440 544948
rect 13 544268 583586 544548
rect 560 543868 583586 544268
rect 13 540868 583586 543868
rect 13 540468 583440 540868
rect 13 540188 583586 540468
rect 560 539788 583586 540188
rect 13 536788 583586 539788
rect 560 536388 583440 536788
rect 13 532708 583586 536388
rect 560 532308 583440 532708
rect 13 528628 583586 532308
rect 560 528228 583440 528628
rect 13 524548 583586 528228
rect 560 524148 583440 524548
rect 13 521148 583586 524148
rect 13 520748 583440 521148
rect 13 520468 583586 520748
rect 560 520068 583586 520468
rect 13 517068 583586 520068
rect 13 516668 583440 517068
rect 13 516388 583586 516668
rect 560 515988 583586 516388
rect 13 512988 583586 515988
rect 13 512588 583440 512988
rect 13 512308 583586 512588
rect 560 511908 583586 512308
rect 13 508908 583586 511908
rect 13 508508 583440 508908
rect 13 508228 583586 508508
rect 560 507828 583586 508228
rect 13 504828 583586 507828
rect 13 504428 583440 504828
rect 13 504148 583586 504428
rect 560 503748 583586 504148
rect 13 500748 583586 503748
rect 13 500348 583440 500748
rect 13 500068 583586 500348
rect 560 499668 583586 500068
rect 13 496668 583586 499668
rect 13 496268 583440 496668
rect 13 495988 583586 496268
rect 560 495588 583586 495988
rect 13 492588 583586 495588
rect 13 492188 583440 492588
rect 13 491908 583586 492188
rect 560 491508 583586 491908
rect 13 488508 583586 491508
rect 13 488108 583440 488508
rect 13 487828 583586 488108
rect 560 487428 583586 487828
rect 13 484428 583586 487428
rect 13 484028 583440 484428
rect 13 483748 583586 484028
rect 560 483348 583586 483748
rect 13 480348 583586 483348
rect 560 479948 583440 480348
rect 13 476268 583586 479948
rect 560 475868 583440 476268
rect 13 472188 583586 475868
rect 560 471788 583440 472188
rect 13 468108 583586 471788
rect 560 467708 583440 468108
rect 13 464028 583586 467708
rect 560 463628 583440 464028
rect 13 460628 583586 463628
rect 13 460228 583440 460628
rect 13 459948 583586 460228
rect 560 459548 583586 459948
rect 13 456548 583586 459548
rect 13 456148 583440 456548
rect 13 455868 583586 456148
rect 560 455468 583586 455868
rect 13 452468 583586 455468
rect 13 452068 583440 452468
rect 13 451788 583586 452068
rect 560 451388 583586 451788
rect 13 448388 583586 451388
rect 13 447988 583440 448388
rect 13 447708 583586 447988
rect 560 447308 583586 447708
rect 13 444308 583586 447308
rect 13 443908 583440 444308
rect 13 443628 583586 443908
rect 560 443228 583586 443628
rect 13 440228 583586 443228
rect 13 439828 583440 440228
rect 13 439548 583586 439828
rect 560 439148 583586 439548
rect 13 436148 583586 439148
rect 13 435748 583440 436148
rect 13 435468 583586 435748
rect 560 435068 583586 435468
rect 13 432068 583586 435068
rect 13 431668 583440 432068
rect 13 431388 583586 431668
rect 560 430988 583586 431388
rect 13 427988 583586 430988
rect 13 427588 583440 427988
rect 13 427308 583586 427588
rect 560 426908 583586 427308
rect 13 423908 583586 426908
rect 13 423508 583440 423908
rect 13 423228 583586 423508
rect 560 422828 583586 423228
rect 13 419828 583586 422828
rect 560 419428 583440 419828
rect 13 415748 583586 419428
rect 560 415348 583440 415748
rect 13 411668 583586 415348
rect 560 411268 583440 411668
rect 13 407588 583586 411268
rect 560 407188 583440 407588
rect 13 404188 583586 407188
rect 13 403788 583440 404188
rect 13 403508 583586 403788
rect 560 403108 583586 403508
rect 13 400108 583586 403108
rect 13 399708 583440 400108
rect 13 399428 583586 399708
rect 560 399028 583586 399428
rect 13 396028 583586 399028
rect 13 395628 583440 396028
rect 13 395348 583586 395628
rect 560 394948 583586 395348
rect 13 391948 583586 394948
rect 13 391548 583440 391948
rect 13 391268 583586 391548
rect 560 390868 583586 391268
rect 13 387868 583586 390868
rect 13 387468 583440 387868
rect 13 387188 583586 387468
rect 560 386788 583586 387188
rect 13 383788 583586 386788
rect 13 383388 583440 383788
rect 13 383108 583586 383388
rect 560 382708 583586 383108
rect 13 379708 583586 382708
rect 13 379308 583440 379708
rect 13 379028 583586 379308
rect 560 378628 583586 379028
rect 13 375628 583586 378628
rect 13 375228 583440 375628
rect 13 374948 583586 375228
rect 560 374548 583586 374948
rect 13 371548 583586 374548
rect 13 371148 583440 371548
rect 13 370868 583586 371148
rect 560 370468 583586 370868
rect 13 367468 583586 370468
rect 13 367068 583440 367468
rect 13 366788 583586 367068
rect 560 366388 583586 366788
rect 13 363388 583586 366388
rect 13 362988 583440 363388
rect 13 362708 583586 362988
rect 560 362308 583586 362708
rect 13 359308 583586 362308
rect 560 358908 583440 359308
rect 13 355228 583586 358908
rect 560 354828 583440 355228
rect 13 351148 583586 354828
rect 560 350748 583440 351148
rect 13 347068 583586 350748
rect 560 346668 583440 347068
rect 13 343668 583586 346668
rect 13 343268 583440 343668
rect 13 342988 583586 343268
rect 560 342588 583586 342988
rect 13 339588 583586 342588
rect 13 339188 583440 339588
rect 13 338908 583586 339188
rect 560 338508 583586 338908
rect 13 335508 583586 338508
rect 13 335108 583440 335508
rect 13 334828 583586 335108
rect 560 334428 583586 334828
rect 13 331428 583586 334428
rect 13 331028 583440 331428
rect 13 330748 583586 331028
rect 560 330348 583586 330748
rect 13 327348 583586 330348
rect 13 326948 583440 327348
rect 13 326668 583586 326948
rect 560 326268 583586 326668
rect 13 323268 583586 326268
rect 13 322868 583440 323268
rect 13 322588 583586 322868
rect 560 322188 583586 322588
rect 13 319188 583586 322188
rect 13 318788 583440 319188
rect 13 318508 583586 318788
rect 560 318108 583586 318508
rect 13 315108 583586 318108
rect 13 314708 583440 315108
rect 13 314428 583586 314708
rect 560 314028 583586 314428
rect 13 311028 583586 314028
rect 13 310628 583440 311028
rect 13 310348 583586 310628
rect 560 309948 583586 310348
rect 13 306948 583586 309948
rect 13 306548 583440 306948
rect 13 306268 583586 306548
rect 560 305868 583586 306268
rect 13 302868 583586 305868
rect 13 302468 583440 302868
rect 13 302188 583586 302468
rect 560 301788 583586 302188
rect 13 298788 583586 301788
rect 560 298388 583440 298788
rect 13 294708 583586 298388
rect 560 294308 583440 294708
rect 13 290628 583586 294308
rect 560 290228 583440 290628
rect 13 286548 583586 290228
rect 560 286148 583440 286548
rect 13 283148 583586 286148
rect 13 282748 583440 283148
rect 13 282468 583586 282748
rect 560 282068 583586 282468
rect 13 279068 583586 282068
rect 13 278668 583440 279068
rect 13 278388 583586 278668
rect 560 277988 583586 278388
rect 13 274988 583586 277988
rect 13 274588 583440 274988
rect 13 274308 583586 274588
rect 560 273908 583586 274308
rect 13 270908 583586 273908
rect 13 270508 583440 270908
rect 13 270228 583586 270508
rect 560 269828 583586 270228
rect 13 266828 583586 269828
rect 13 266428 583440 266828
rect 13 266148 583586 266428
rect 560 265748 583586 266148
rect 13 262748 583586 265748
rect 13 262348 583440 262748
rect 13 262068 583586 262348
rect 560 261668 583586 262068
rect 13 258668 583586 261668
rect 13 258268 583440 258668
rect 13 257988 583586 258268
rect 560 257588 583586 257988
rect 13 254588 583586 257588
rect 13 254188 583440 254588
rect 13 253908 583586 254188
rect 560 253508 583586 253908
rect 13 250508 583586 253508
rect 13 250108 583440 250508
rect 13 249828 583586 250108
rect 560 249428 583586 249828
rect 13 246428 583586 249428
rect 13 246028 583440 246428
rect 13 245748 583586 246028
rect 560 245348 583586 245748
rect 13 242348 583586 245348
rect 13 241948 583440 242348
rect 13 241668 583586 241948
rect 560 241268 583586 241668
rect 13 238268 583586 241268
rect 560 237868 583440 238268
rect 13 234188 583586 237868
rect 560 233788 583440 234188
rect 13 230108 583586 233788
rect 560 229708 583440 230108
rect 13 226028 583586 229708
rect 560 225628 583440 226028
rect 13 222628 583586 225628
rect 13 222228 583440 222628
rect 13 221948 583586 222228
rect 560 221548 583586 221948
rect 13 218548 583586 221548
rect 13 218148 583440 218548
rect 13 217868 583586 218148
rect 560 217468 583586 217868
rect 13 214468 583586 217468
rect 13 214068 583440 214468
rect 13 213788 583586 214068
rect 560 213388 583586 213788
rect 13 210388 583586 213388
rect 13 209988 583440 210388
rect 13 209708 583586 209988
rect 560 209308 583586 209708
rect 13 206308 583586 209308
rect 13 205908 583440 206308
rect 13 205628 583586 205908
rect 560 205228 583586 205628
rect 13 202228 583586 205228
rect 13 201828 583440 202228
rect 13 201548 583586 201828
rect 560 201148 583586 201548
rect 13 198148 583586 201148
rect 13 197748 583440 198148
rect 13 197468 583586 197748
rect 560 197068 583586 197468
rect 13 194068 583586 197068
rect 13 193668 583440 194068
rect 13 193388 583586 193668
rect 560 192988 583586 193388
rect 13 189988 583586 192988
rect 13 189588 583440 189988
rect 13 189308 583586 189588
rect 560 188908 583586 189308
rect 13 185908 583586 188908
rect 13 185508 583440 185908
rect 13 185228 583586 185508
rect 560 184828 583586 185228
rect 13 181828 583586 184828
rect 13 181428 583440 181828
rect 13 181148 583586 181428
rect 560 180748 583586 181148
rect 13 177748 583586 180748
rect 560 177348 583440 177748
rect 13 173668 583586 177348
rect 560 173268 583440 173668
rect 13 169588 583586 173268
rect 560 169188 583440 169588
rect 13 165508 583586 169188
rect 560 165108 583440 165508
rect 13 162108 583586 165108
rect 13 161708 583440 162108
rect 13 161428 583586 161708
rect 560 161028 583586 161428
rect 13 158028 583586 161028
rect 13 157628 583440 158028
rect 13 157348 583586 157628
rect 560 156948 583586 157348
rect 13 153948 583586 156948
rect 13 153548 583440 153948
rect 13 153268 583586 153548
rect 560 152868 583586 153268
rect 13 149868 583586 152868
rect 13 149468 583440 149868
rect 13 149188 583586 149468
rect 560 148788 583586 149188
rect 13 145788 583586 148788
rect 13 145388 583440 145788
rect 13 145108 583586 145388
rect 560 144708 583586 145108
rect 13 141708 583586 144708
rect 13 141308 583440 141708
rect 13 141028 583586 141308
rect 560 140628 583586 141028
rect 13 137628 583586 140628
rect 13 137228 583440 137628
rect 13 136948 583586 137228
rect 560 136548 583586 136948
rect 13 133548 583586 136548
rect 13 133148 583440 133548
rect 13 132868 583586 133148
rect 560 132468 583586 132868
rect 13 129468 583586 132468
rect 13 129068 583440 129468
rect 13 128788 583586 129068
rect 560 128388 583586 128788
rect 13 125388 583586 128388
rect 13 124988 583440 125388
rect 13 124708 583586 124988
rect 560 124308 583586 124708
rect 13 121308 583586 124308
rect 13 120908 583440 121308
rect 13 120628 583586 120908
rect 560 120228 583586 120628
rect 13 117228 583586 120228
rect 560 116828 583440 117228
rect 13 113148 583586 116828
rect 560 112748 583440 113148
rect 13 109068 583586 112748
rect 560 108668 583440 109068
rect 13 104988 583586 108668
rect 560 104588 583440 104988
rect 13 101588 583586 104588
rect 13 101188 583440 101588
rect 13 100908 583586 101188
rect 560 100508 583586 100908
rect 13 97508 583586 100508
rect 13 97108 583440 97508
rect 13 96828 583586 97108
rect 560 96428 583586 96828
rect 13 93428 583586 96428
rect 13 93028 583440 93428
rect 13 92748 583586 93028
rect 560 92348 583586 92748
rect 13 89348 583586 92348
rect 13 88948 583440 89348
rect 13 88668 583586 88948
rect 560 88268 583586 88668
rect 13 85268 583586 88268
rect 13 84868 583440 85268
rect 13 84588 583586 84868
rect 560 84188 583586 84588
rect 13 81188 583586 84188
rect 13 80788 583440 81188
rect 13 80508 583586 80788
rect 560 80108 583586 80508
rect 13 77108 583586 80108
rect 13 76708 583440 77108
rect 13 76428 583586 76708
rect 560 76028 583586 76428
rect 13 73028 583586 76028
rect 13 72628 583440 73028
rect 13 72348 583586 72628
rect 560 71948 583586 72348
rect 13 68948 583586 71948
rect 13 68548 583440 68948
rect 13 68268 583586 68548
rect 560 67868 583586 68268
rect 13 64868 583586 67868
rect 13 64468 583440 64868
rect 13 64188 583586 64468
rect 560 63788 583586 64188
rect 13 60788 583586 63788
rect 13 60388 583440 60788
rect 13 60108 583586 60388
rect 560 59708 583586 60108
rect 13 56708 583586 59708
rect 560 56308 583440 56708
rect 13 52628 583586 56308
rect 560 52228 583440 52628
rect 13 48548 583586 52228
rect 560 48148 583440 48548
rect 13 44468 583586 48148
rect 560 44068 583440 44468
rect 13 41068 583586 44068
rect 13 40668 583440 41068
rect 13 40388 583586 40668
rect 560 39988 583586 40388
rect 13 36988 583586 39988
rect 13 36588 583440 36988
rect 13 36308 583586 36588
rect 560 35908 583586 36308
rect 13 32908 583586 35908
rect 13 32508 583440 32908
rect 13 32228 583586 32508
rect 560 31828 583586 32228
rect 13 28828 583586 31828
rect 13 28428 583440 28828
rect 13 28148 583586 28428
rect 560 27748 583586 28148
rect 13 24748 583586 27748
rect 13 24348 583440 24748
rect 13 24068 583586 24348
rect 560 23668 583586 24068
rect 13 20668 583586 23668
rect 13 20268 583440 20668
rect 13 19988 583586 20268
rect 560 19588 583586 19988
rect 13 16588 583586 19588
rect 13 16188 583440 16588
rect 13 15908 583586 16188
rect 560 15508 583586 15908
rect 13 12508 583586 15508
rect 13 12108 583440 12508
rect 13 11828 583586 12108
rect 560 11428 583586 11828
rect 13 8428 583586 11428
rect 13 8028 583440 8428
rect 13 7748 583586 8028
rect 560 7348 583586 7748
rect 13 4348 583586 7348
rect 13 3948 583440 4348
rect 13 3668 583586 3948
rect 560 3268 583586 3668
rect 13 268 583586 3268
rect 13 35 583440 268
<< metal4 >>
rect -8726 -7654 -8106 711590
rect -7766 -6694 -7146 710630
rect -6806 -5734 -6186 709670
rect -5846 -4774 -5226 708710
rect -4886 -3814 -4266 707750
rect -3926 -2854 -3306 706790
rect -2966 -1894 -2346 705830
rect -2006 -934 -1386 704870
rect 1794 -7654 2414 711590
rect 5514 -7654 6134 711590
rect 9234 -7654 9854 711590
rect 12954 -7654 13574 711590
rect 16674 -7654 17294 711590
rect 20394 -7654 21014 711590
rect 24114 -7654 24734 711590
rect 27834 -7654 28454 711590
rect 37794 -7654 38414 711590
rect 41514 -7654 42134 711590
rect 45234 -7654 45854 711590
rect 48954 -7654 49574 711590
rect 52674 -7654 53294 711590
rect 56394 -7654 57014 711590
rect 60114 -7654 60734 711590
rect 63834 -7654 64454 711590
rect 73794 -7654 74414 711590
rect 77514 -7654 78134 711590
rect 81234 -7654 81854 711590
rect 84954 -7654 85574 711590
rect 88674 -7654 89294 711590
rect 92394 -7654 93014 711590
rect 96114 -7654 96734 711590
rect 99834 -7654 100454 711590
rect 109794 -7654 110414 711590
rect 113514 -7654 114134 711590
rect 117234 -7654 117854 711590
rect 120954 -7654 121574 711590
rect 124674 -7654 125294 711590
rect 128394 -7654 129014 711590
rect 132114 -7654 132734 711590
rect 135834 -7654 136454 711590
rect 145794 -7654 146414 711590
rect 149514 -7654 150134 711590
rect 153234 -7654 153854 711590
rect 156954 -7654 157574 711590
rect 160674 -7654 161294 711590
rect 164394 -7654 165014 711590
rect 168114 -7654 168734 711590
rect 171834 -7654 172454 711590
rect 181794 -7654 182414 711590
rect 185514 -7654 186134 711590
rect 189234 -7654 189854 711590
rect 192954 -7654 193574 711590
rect 196674 -7654 197294 711590
rect 200394 -7654 201014 711590
rect 204114 -7654 204734 711590
rect 207834 -7654 208454 711590
rect 217794 -7654 218414 711590
rect 221514 -7654 222134 711590
rect 225234 -7654 225854 711590
rect 228954 -7654 229574 711590
rect 232674 -7654 233294 711590
rect 236394 -7654 237014 711590
rect 240114 -7654 240734 711590
rect 243834 -7654 244454 711590
rect 253794 -7654 254414 711590
rect 257514 -7654 258134 711590
rect 261234 -7654 261854 711590
rect 264954 -7654 265574 711590
rect 268674 -7654 269294 711590
rect 272394 -7654 273014 711590
rect 276114 -7654 276734 711590
rect 279834 -7654 280454 711590
rect 289794 -7654 290414 711590
rect 293514 -7654 294134 711590
rect 297234 -7654 297854 711590
rect 300954 -7654 301574 711590
rect 304674 -7654 305294 711590
rect 308394 -7654 309014 711590
rect 312114 -7654 312734 711590
rect 315834 -7654 316454 711590
rect 325794 -7654 326414 711590
rect 329514 -7654 330134 711590
rect 333234 -7654 333854 711590
rect 336954 -7654 337574 711590
rect 340674 -7654 341294 711590
rect 344394 -7654 345014 711590
rect 348114 -7654 348734 711590
rect 351834 -7654 352454 711590
rect 361794 -7654 362414 711590
rect 365514 -7654 366134 711590
rect 369234 -7654 369854 711590
rect 372954 -7654 373574 711590
rect 376674 -7654 377294 711590
rect 380394 -7654 381014 711590
rect 384114 -7654 384734 711590
rect 387834 -7654 388454 711590
rect 397794 -7654 398414 711590
rect 401514 -7654 402134 711590
rect 405234 -7654 405854 711590
rect 408954 -7654 409574 711590
rect 412674 -7654 413294 711590
rect 416394 -7654 417014 711590
rect 420114 -7654 420734 711590
rect 423834 -7654 424454 711590
rect 433794 -7654 434414 711590
rect 437514 -7654 438134 711590
rect 441234 -7654 441854 711590
rect 444954 -7654 445574 711590
rect 448674 -7654 449294 711590
rect 452394 -7654 453014 711590
rect 456114 -7654 456734 711590
rect 459834 -7654 460454 711590
rect 469794 -7654 470414 711590
rect 473514 -7654 474134 711590
rect 477234 -7654 477854 711590
rect 480954 -7654 481574 711590
rect 484674 -7654 485294 711590
rect 488394 -7654 489014 711590
rect 492114 -7654 492734 711590
rect 495834 -7654 496454 711590
rect 505794 -7654 506414 711590
rect 509514 -7654 510134 711590
rect 513234 -7654 513854 711590
rect 516954 -7654 517574 711590
rect 520674 -7654 521294 711590
rect 524394 -7654 525014 711590
rect 528114 -7654 528734 711590
rect 531834 -7654 532454 711590
rect 541794 -7654 542414 711590
rect 545514 -7654 546134 711590
rect 549234 -7654 549854 711590
rect 552954 -7654 553574 711590
rect 556674 -7654 557294 711590
rect 560394 -7654 561014 711590
rect 564114 -7654 564734 711590
rect 567834 -7654 568454 711590
rect 577794 -7654 578414 711590
rect 581514 -7654 582134 711590
rect 585310 -934 585930 704870
rect 586270 -1894 586890 705830
rect 587230 -2854 587850 706790
rect 588190 -3814 588810 707750
rect 589150 -4774 589770 708710
rect 590110 -5734 590730 709670
rect 591070 -6694 591690 710630
rect 592030 -7654 592650 711590
<< obsm4 >>
rect 3187 3299 5434 699821
rect 6214 3299 9154 699821
rect 9934 3299 12874 699821
rect 13654 3299 16594 699821
rect 17374 3299 20314 699821
rect 21094 3299 24034 699821
rect 24814 3299 27754 699821
rect 28534 3299 37714 699821
rect 38494 3299 41434 699821
rect 42214 3299 45154 699821
rect 45934 3299 48874 699821
rect 49654 3299 52594 699821
rect 53374 3299 56314 699821
rect 57094 3299 60034 699821
rect 60814 3299 63754 699821
rect 64534 3299 73714 699821
rect 74494 3299 77434 699821
rect 78214 3299 81154 699821
rect 81934 3299 84874 699821
rect 85654 3299 88594 699821
rect 89374 3299 92314 699821
rect 93094 3299 96034 699821
rect 96814 3299 99754 699821
rect 100534 3299 109714 699821
rect 110494 3299 113434 699821
rect 114214 3299 117154 699821
rect 117934 3299 120874 699821
rect 121654 3299 124594 699821
rect 125374 3299 128314 699821
rect 129094 3299 132034 699821
rect 132814 3299 135754 699821
rect 136534 3299 145714 699821
rect 146494 3299 149434 699821
rect 150214 3299 153154 699821
rect 153934 3299 156874 699821
rect 157654 3299 160594 699821
rect 161374 3299 164314 699821
rect 165094 3299 168034 699821
rect 168814 3299 171754 699821
rect 172534 3299 181714 699821
rect 182494 3299 185434 699821
rect 186214 3299 189154 699821
rect 189934 3299 192874 699821
rect 193654 3299 196594 699821
rect 197374 3299 200314 699821
rect 201094 3299 204034 699821
rect 204814 3299 207754 699821
rect 208534 3299 217714 699821
rect 218494 3299 221434 699821
rect 222214 3299 225154 699821
rect 225934 3299 228874 699821
rect 229654 3299 232594 699821
rect 233374 3299 236314 699821
rect 237094 3299 240034 699821
rect 240814 3299 243754 699821
rect 244534 3299 253714 699821
rect 254494 3299 257434 699821
rect 258214 3299 261154 699821
rect 261934 3299 264874 699821
rect 265654 3299 268594 699821
rect 269374 3299 272314 699821
rect 273094 3299 276034 699821
rect 276814 3299 279754 699821
rect 280534 3299 289714 699821
rect 290494 3299 293434 699821
rect 294214 3299 297154 699821
rect 297934 3299 300874 699821
rect 301654 3299 304594 699821
rect 305374 3299 308314 699821
rect 309094 3299 312034 699821
rect 312814 3299 315754 699821
rect 316534 3299 325714 699821
rect 326494 3299 329434 699821
rect 330214 3299 333154 699821
rect 333934 3299 336874 699821
rect 337654 3299 340594 699821
rect 341374 3299 344314 699821
rect 345094 3299 348034 699821
rect 348814 3299 351754 699821
rect 352534 3299 361714 699821
rect 362494 3299 365434 699821
rect 366214 3299 369154 699821
rect 369934 3299 372874 699821
rect 373654 3299 376594 699821
rect 377374 3299 380314 699821
rect 381094 3299 384034 699821
rect 384814 3299 387754 699821
rect 388534 3299 397714 699821
rect 398494 3299 401434 699821
rect 402214 3299 405154 699821
rect 405934 3299 408874 699821
rect 409654 3299 412594 699821
rect 413374 3299 416314 699821
rect 417094 3299 420034 699821
rect 420814 3299 423754 699821
rect 424534 3299 433714 699821
rect 434494 3299 437434 699821
rect 438214 3299 441154 699821
rect 441934 3299 444874 699821
rect 445654 3299 448594 699821
rect 449374 3299 452314 699821
rect 453094 3299 456034 699821
rect 456814 3299 459754 699821
rect 460534 3299 469714 699821
rect 470494 3299 473434 699821
rect 474214 3299 477154 699821
rect 477934 3299 480874 699821
rect 481654 3299 484594 699821
rect 485374 3299 488314 699821
rect 489094 3299 492034 699821
rect 492814 3299 495754 699821
rect 496534 3299 505714 699821
rect 506494 3299 509434 699821
rect 510214 3299 513154 699821
rect 513934 3299 516874 699821
rect 517654 3299 520594 699821
rect 521374 3299 524314 699821
rect 525094 3299 528034 699821
rect 528814 3299 531754 699821
rect 532534 3299 541714 699821
rect 542494 3299 545434 699821
rect 546214 3299 549154 699821
rect 549934 3299 552874 699821
rect 553654 3299 556594 699821
rect 557374 3299 560314 699821
rect 561094 3299 564034 699821
rect 564814 3299 567754 699821
rect 568534 3299 577714 699821
rect 578494 3299 581197 699821
<< metal5 >>
rect -8726 710970 592650 711590
rect -7766 710010 591690 710630
rect -6806 709050 590730 709670
rect -5846 708090 589770 708710
rect -4886 707130 588810 707750
rect -3926 706170 587850 706790
rect -2966 705210 586890 705830
rect -2006 704250 585930 704870
rect -8726 698026 592650 698646
rect -8726 694306 592650 694926
rect -8726 690586 592650 691206
rect -8726 686866 592650 687486
rect -8726 676906 592650 677526
rect -8726 673186 592650 673806
rect -8726 669466 592650 670086
rect -8726 665746 592650 666366
rect -8726 662026 592650 662646
rect -8726 658306 592650 658926
rect -8726 654586 592650 655206
rect -8726 650866 592650 651486
rect -8726 640906 592650 641526
rect -8726 637186 592650 637806
rect -8726 633466 592650 634086
rect -8726 629746 592650 630366
rect -8726 626026 592650 626646
rect -8726 622306 592650 622926
rect -8726 618586 592650 619206
rect -8726 614866 592650 615486
rect -8726 604906 592650 605526
rect -8726 601186 592650 601806
rect -8726 597466 592650 598086
rect -8726 593746 592650 594366
rect -8726 590026 592650 590646
rect -8726 586306 592650 586926
rect -8726 582586 592650 583206
rect -8726 578866 592650 579486
rect -8726 568906 592650 569526
rect -8726 565186 592650 565806
rect -8726 561466 592650 562086
rect -8726 557746 592650 558366
rect -8726 554026 592650 554646
rect -8726 550306 592650 550926
rect -8726 546586 592650 547206
rect -8726 542866 592650 543486
rect -8726 532906 592650 533526
rect -8726 529186 592650 529806
rect -8726 525466 592650 526086
rect -8726 521746 592650 522366
rect -8726 518026 592650 518646
rect -8726 514306 592650 514926
rect -8726 510586 592650 511206
rect -8726 506866 592650 507486
rect -8726 496906 592650 497526
rect -8726 493186 592650 493806
rect -8726 489466 592650 490086
rect -8726 485746 592650 486366
rect -8726 482026 592650 482646
rect -8726 478306 592650 478926
rect -8726 474586 592650 475206
rect -8726 470866 592650 471486
rect -8726 460906 592650 461526
rect -8726 457186 592650 457806
rect -8726 453466 592650 454086
rect -8726 449746 592650 450366
rect -8726 446026 592650 446646
rect -8726 442306 592650 442926
rect -8726 438586 592650 439206
rect -8726 434866 592650 435486
rect -8726 424906 592650 425526
rect -8726 421186 592650 421806
rect -8726 417466 592650 418086
rect -8726 413746 592650 414366
rect -8726 410026 592650 410646
rect -8726 406306 592650 406926
rect -8726 402586 592650 403206
rect -8726 398866 592650 399486
rect -8726 388906 592650 389526
rect -8726 385186 592650 385806
rect -8726 381466 592650 382086
rect -8726 377746 592650 378366
rect -8726 374026 592650 374646
rect -8726 370306 592650 370926
rect -8726 366586 592650 367206
rect -8726 362866 592650 363486
rect -8726 352906 592650 353526
rect -8726 349186 592650 349806
rect -8726 345466 592650 346086
rect -8726 341746 592650 342366
rect -8726 338026 592650 338646
rect -8726 334306 592650 334926
rect -8726 330586 592650 331206
rect -8726 326866 592650 327486
rect -8726 316906 592650 317526
rect -8726 313186 592650 313806
rect -8726 309466 592650 310086
rect -8726 305746 592650 306366
rect -8726 302026 592650 302646
rect -8726 298306 592650 298926
rect -8726 294586 592650 295206
rect -8726 290866 592650 291486
rect -8726 280906 592650 281526
rect -8726 277186 592650 277806
rect -8726 273466 592650 274086
rect -8726 269746 592650 270366
rect -8726 266026 592650 266646
rect -8726 262306 592650 262926
rect -8726 258586 592650 259206
rect -8726 254866 592650 255486
rect -8726 244906 592650 245526
rect -8726 241186 592650 241806
rect -8726 237466 592650 238086
rect -8726 233746 592650 234366
rect -8726 230026 592650 230646
rect -8726 226306 592650 226926
rect -8726 222586 592650 223206
rect -8726 218866 592650 219486
rect -8726 208906 592650 209526
rect -8726 205186 592650 205806
rect -8726 201466 592650 202086
rect -8726 197746 592650 198366
rect -8726 194026 592650 194646
rect -8726 190306 592650 190926
rect -8726 186586 592650 187206
rect -8726 182866 592650 183486
rect -8726 172906 592650 173526
rect -8726 169186 592650 169806
rect -8726 165466 592650 166086
rect -8726 161746 592650 162366
rect -8726 158026 592650 158646
rect -8726 154306 592650 154926
rect -8726 150586 592650 151206
rect -8726 146866 592650 147486
rect -8726 136906 592650 137526
rect -8726 133186 592650 133806
rect -8726 129466 592650 130086
rect -8726 125746 592650 126366
rect -8726 122026 592650 122646
rect -8726 118306 592650 118926
rect -8726 114586 592650 115206
rect -8726 110866 592650 111486
rect -8726 100906 592650 101526
rect -8726 97186 592650 97806
rect -8726 93466 592650 94086
rect -8726 89746 592650 90366
rect -8726 86026 592650 86646
rect -8726 82306 592650 82926
rect -8726 78586 592650 79206
rect -8726 74866 592650 75486
rect -8726 64906 592650 65526
rect -8726 61186 592650 61806
rect -8726 57466 592650 58086
rect -8726 53746 592650 54366
rect -8726 50026 592650 50646
rect -8726 46306 592650 46926
rect -8726 42586 592650 43206
rect -8726 38866 592650 39486
rect -8726 28906 592650 29526
rect -8726 25186 592650 25806
rect -8726 21466 592650 22086
rect -8726 17746 592650 18366
rect -8726 14026 592650 14646
rect -8726 10306 592650 10926
rect -8726 6586 592650 7206
rect -8726 2866 592650 3486
rect -2006 -934 585930 -314
rect -2966 -1894 586890 -1274
rect -3926 -2854 587850 -2234
rect -4886 -3814 588810 -3194
rect -5846 -4774 589770 -4154
rect -6806 -5734 590730 -5114
rect -7766 -6694 591690 -6074
rect -8726 -7654 592650 -7034
<< labels >>
rlabel metal2 s 87574 -960 87686 480 8 gpio_analog[0]
port 1 nsew
rlabel metal2 s 156482 -960 156594 480 8 gpio_analog[10]
port 2 nsew
rlabel metal3 s 583520 56388 584960 56628 6 gpio_analog[11]
port 3 nsew
rlabel metal2 s 100454 703520 100566 704960 6 gpio_analog[12]
port 4 nsew
rlabel metal3 s -960 326348 480 326588 4 gpio_analog[13]
port 5 nsew
rlabel metal2 s 345174 703520 345286 704960 6 gpio_analog[14]
port 6 nsew
rlabel metal3 s 583520 222308 584960 222548 6 gpio_analog[15]
port 7 nsew
rlabel metal3 s -960 637108 480 637348 4 gpio_analog[16]
port 8 nsew
rlabel metal3 s -960 128468 480 128708 4 gpio_analog[17]
port 9 nsew
rlabel metal3 s 583520 80868 584960 81108 6 gpio_analog[1]
port 10 nsew
rlabel metal2 s 259522 -960 259634 480 8 gpio_analog[2]
port 11 nsew
rlabel metal3 s -960 435148 480 435388 4 gpio_analog[3]
port 12 nsew
rlabel metal3 s 583520 673828 584960 674068 6 gpio_analog[4]
port 13 nsew
rlabel metal3 s -960 205308 480 205548 4 gpio_analog[5]
port 14 nsew
rlabel metal3 s -960 399108 480 399348 4 gpio_analog[6]
port 15 nsew
rlabel metal2 s 75982 -960 76094 480 8 gpio_analog[7]
port 16 nsew
rlabel metal2 s 546102 -960 546214 480 8 gpio_analog[8]
port 17 nsew
rlabel metal2 s 412150 -960 412262 480 8 gpio_analog[9]
port 18 nsew
rlabel metal2 s 240202 -960 240314 480 8 gpio_noesd[0]
port 19 nsew
rlabel metal3 s -960 536468 480 536708 4 gpio_noesd[10]
port 20 nsew
rlabel metal3 s -960 447388 480 447628 4 gpio_noesd[11]
port 21 nsew
rlabel metal2 s 173226 703520 173338 704960 6 gpio_noesd[12]
port 22 nsew
rlabel metal2 s 390898 703520 391010 704960 6 gpio_noesd[13]
port 23 nsew
rlabel metal3 s -960 382788 480 383028 4 gpio_noesd[14]
port 24 nsew
rlabel metal3 s -960 59788 480 60028 4 gpio_noesd[15]
port 25 nsew
rlabel metal3 s 583520 28508 584960 28748 6 gpio_noesd[16]
port 26 nsew
rlabel metal2 s 211222 703520 211334 704960 6 gpio_noesd[17]
port 27 nsew
rlabel metal2 s 121706 -960 121818 480 8 gpio_noesd[1]
port 28 nsew
rlabel metal2 s 328430 -960 328542 480 8 gpio_noesd[2]
port 29 nsew
rlabel metal3 s 583520 641868 584960 642108 6 gpio_noesd[3]
port 30 nsew
rlabel metal2 s 191902 703520 192014 704960 6 gpio_noesd[4]
port 31 nsew
rlabel metal3 s 583520 64548 584960 64788 6 gpio_noesd[5]
port 32 nsew
rlabel metal3 s 583520 601068 584960 601308 6 gpio_noesd[6]
port 33 nsew
rlabel metal3 s 583520 492268 584960 492508 6 gpio_noesd[7]
port 34 nsew
rlabel metal3 s -960 88348 480 88588 4 gpio_noesd[8]
port 35 nsew
rlabel metal3 s -960 132548 480 132788 4 gpio_noesd[9]
port 36 nsew
rlabel metal3 s -960 245428 480 245668 4 io_analog[0]
port 37 nsew
rlabel metal2 s 56662 -960 56774 480 8 io_analog[10]
port 38 nsew
rlabel metal3 s 583520 60468 584960 60708 6 io_analog[1]
port 39 nsew
rlabel metal3 s 583520 552788 584960 553028 6 io_analog[2]
port 40 nsew
rlabel metal2 s 228610 -960 228722 480 8 io_analog[3]
port 41 nsew
rlabel metal2 s 113978 -960 114090 480 8 io_analog[4]
port 42 nsew
rlabel metal2 s 88862 703520 88974 704960 6 io_analog[5]
port 43 nsew
rlabel metal2 s 450790 -960 450902 480 8 io_analog[6]
port 44 nsew
rlabel metal3 s -960 233868 480 234108 4 io_analog[7]
port 45 nsew
rlabel metal2 s 209934 -960 210046 480 8 io_analog[8]
port 46 nsew
rlabel metal3 s -960 334508 480 334748 4 io_analog[9]
port 47 nsew
rlabel metal2 s 22530 -960 22642 480 8 io_clamp_high[0]
port 48 nsew
rlabel metal3 s 583520 581348 584960 581588 6 io_clamp_high[1]
port 49 nsew
rlabel metal3 s 583520 363068 584960 363308 6 io_clamp_high[2]
port 50 nsew
rlabel metal3 s -960 124388 480 124628 4 io_clamp_low[0]
port 51 nsew
rlabel metal2 s 285926 -960 286038 480 8 io_clamp_low[1]
port 52 nsew
rlabel metal3 s -960 649348 480 649588 4 io_clamp_low[2]
port 53 nsew
rlabel metal2 s 37986 -960 38098 480 8 io_in[0]
port 54 nsew
rlabel metal3 s 583520 504508 584960 504748 6 io_in[10]
port 55 nsew
rlabel metal2 s 493938 703520 494050 704960 6 io_in[11]
port 56 nsew
rlabel metal2 s 402490 703520 402602 704960 6 io_in[12]
port 57 nsew
rlabel metal2 s 99166 -960 99278 480 8 io_in[13]
port 58 nsew
rlabel metal2 s 416014 -960 416126 480 8 io_in[14]
port 59 nsew
rlabel metal3 s -960 76108 480 76348 4 io_in[15]
port 60 nsew
rlabel metal2 s 519054 -960 519166 480 8 io_in[16]
port 61 nsew
rlabel metal3 s 583520 237948 584960 238188 6 io_in[17]
port 62 nsew
rlabel metal3 s 583520 72708 584960 72948 6 io_in[18]
port 63 nsew
rlabel metal3 s -960 564348 480 564588 4 io_in[19]
port 64 nsew
rlabel metal2 s 492650 -960 492762 480 8 io_in[1]
port 65 nsew
rlabel metal2 s 534510 -960 534622 480 8 io_in[20]
port 66 nsew
rlabel metal2 s 336158 -960 336270 480 8 io_in[21]
port 67 nsew
rlabel metal3 s 583520 133228 584960 133468 6 io_in[22]
port 68 nsew
rlabel metal2 s 264674 703520 264786 704960 6 io_in[23]
port 69 nsew
rlabel metal3 s 583520 399788 584960 400028 6 io_in[24]
port 70 nsew
rlabel metal2 s 580234 -960 580346 480 8 io_in[25]
port 71 nsew
rlabel metal2 s 535798 703520 535910 704960 6 io_in[26]
port 72 nsew
rlabel metal3 s 583520 452148 584960 452388 6 io_in[2]
port 73 nsew
rlabel metal3 s -960 314108 480 314348 4 io_in[3]
port 74 nsew
rlabel metal2 s 427606 -960 427718 480 8 io_in[4]
port 75 nsew
rlabel metal2 s 130722 703520 130834 704960 6 io_in[5]
port 76 nsew
rlabel metal3 s 583520 548708 584960 548948 6 io_in[6]
port 77 nsew
rlabel metal3 s -960 56388 480 56628 4 io_in[7]
port 78 nsew
rlabel metal2 s 83710 -960 83822 480 8 io_in[8]
port 79 nsew
rlabel metal2 s 230542 703520 230654 704960 6 io_in[9]
port 80 nsew
rlabel metal2 s 164210 -960 164322 480 8 io_in_3v3[0]
port 81 nsew
rlabel metal2 s 45714 -960 45826 480 8 io_in_3v3[10]
port 82 nsew
rlabel metal2 s 337446 703520 337558 704960 6 io_in_3v3[11]
port 83 nsew
rlabel metal2 s 531934 703520 532046 704960 6 io_in_3v3[12]
port 84 nsew
rlabel metal2 s 10938 -960 11050 480 8 io_in_3v3[13]
port 85 nsew
rlabel metal3 s -960 641188 480 641428 4 io_in_3v3[14]
port 86 nsew
rlabel metal3 s 583520 205988 584960 206228 6 io_in_3v3[15]
port 87 nsew
rlabel metal3 s 583520 157708 584960 157948 6 io_in_3v3[16]
port 88 nsew
rlabel metal3 s -960 657508 480 657748 4 io_in_3v3[17]
port 89 nsew
rlabel metal3 s -960 366468 480 366708 4 io_in_3v3[18]
port 90 nsew
rlabel metal3 s -960 633028 480 633268 4 io_in_3v3[19]
port 91 nsew
rlabel metal3 s 583520 52308 584960 52548 6 io_in_3v3[1]
port 92 nsew
rlabel metal2 s 73406 703520 73518 704960 6 io_in_3v3[20]
port 93 nsew
rlabel metal3 s -960 592908 480 593148 4 io_in_3v3[21]
port 94 nsew
rlabel metal3 s -960 697628 480 697868 4 io_in_3v3[22]
port 95 nsew
rlabel metal3 s -960 677228 480 677468 4 io_in_3v3[23]
port 96 nsew
rlabel metal2 s 293654 -960 293766 480 8 io_in_3v3[24]
port 97 nsew
rlabel metal3 s 583520 335188 584960 335428 6 io_in_3v3[25]
port 98 nsew
rlabel metal3 s -960 395028 480 395268 4 io_in_3v3[26]
port 99 nsew
rlabel metal2 s 1278 703520 1390 704960 6 io_in_3v3[2]
port 100 nsew
rlabel metal3 s 583520 653428 584960 653668 6 io_in_3v3[3]
port 101 nsew
rlabel metal2 s 566710 703520 566822 704960 6 io_in_3v3[4]
port 102 nsew
rlabel metal2 s 312974 -960 313086 480 8 io_in_3v3[5]
port 103 nsew
rlabel metal2 s 446926 -960 447038 480 8 io_in_3v3[6]
port 104 nsew
rlabel metal2 s 198342 -960 198454 480 8 io_in_3v3[7]
port 105 nsew
rlabel metal2 s 295586 703520 295698 704960 6 io_in_3v3[8]
port 106 nsew
rlabel metal2 s 553830 -960 553942 480 8 io_in_3v3[9]
port 107 nsew
rlabel metal3 s -960 475948 480 476188 4 io_oeb[0]
port 108 nsew
rlabel metal2 s 474618 703520 474730 704960 6 io_oeb[10]
port 109 nsew
rlabel metal2 s 218950 703520 219062 704960 6 io_oeb[11]
port 110 nsew
rlabel metal2 s 366426 -960 366538 480 8 io_oeb[12]
port 111 nsew
rlabel metal2 s 515190 -960 515302 480 8 io_oeb[13]
port 112 nsew
rlabel metal3 s 583520 350828 584960 351068 6 io_oeb[14]
port 113 nsew
rlabel metal3 s -960 487508 480 487748 4 io_oeb[15]
port 114 nsew
rlabel metal3 s -960 528308 480 528548 4 io_oeb[16]
port 115 nsew
rlabel metal3 s 583520 592908 584960 593148 6 io_oeb[17]
port 116 nsew
rlabel metal2 s 129434 -960 129546 480 8 io_oeb[18]
port 117 nsew
rlabel metal3 s 583520 649348 584960 649588 6 io_oeb[19]
port 118 nsew
rlabel metal2 s 501666 703520 501778 704960 6 io_oeb[1]
port 119 nsew
rlabel metal2 s 524850 703520 524962 704960 6 io_oeb[20]
port 120 nsew
rlabel metal2 s 478482 703520 478594 704960 6 io_oeb[21]
port 121 nsew
rlabel metal2 s 60526 -960 60638 480 8 io_oeb[22]
port 122 nsew
rlabel metal3 s 583520 169268 584960 169508 6 io_oeb[23]
port 123 nsew
rlabel metal2 s 349038 703520 349150 704960 6 io_oeb[24]
port 124 nsew
rlabel metal3 s 583520 484108 584960 484348 6 io_oeb[25]
port 125 nsew
rlabel metal3 s 583520 375308 584960 375548 6 io_oeb[26]
port 126 nsew
rlabel metal3 s -960 608548 480 608788 4 io_oeb[2]
port 127 nsew
rlabel metal3 s -960 624868 480 625108 4 io_oeb[3]
port 128 nsew
rlabel metal3 s -960 467788 480 468028 4 io_oeb[4]
port 129 nsew
rlabel metal3 s 583520 560948 584960 561188 6 io_oeb[5]
port 130 nsew
rlabel metal2 s 39274 703520 39386 704960 6 io_oeb[6]
port 131 nsew
rlabel metal3 s -960 520148 480 520388 4 io_oeb[7]
port 132 nsew
rlabel metal2 s 299450 703520 299562 704960 6 io_oeb[8]
port 133 nsew
rlabel metal3 s 583520 294388 584960 294628 6 io_oeb[9]
port 134 nsew
rlabel metal2 s 520986 703520 521098 704960 6 io_out[0]
port 135 nsew
rlabel metal3 s -960 177428 480 177668 4 io_out[10]
port 136 nsew
rlabel metal3 s 583520 665668 584960 665908 6 io_out[11]
port 137 nsew
rlabel metal3 s -960 298468 480 298708 4 io_out[12]
port 138 nsew
rlabel metal3 s 583520 415428 584960 415668 6 io_out[13]
port 139 nsew
rlabel metal2 s 268538 703520 268650 704960 6 io_out[14]
port 140 nsew
rlabel metal3 s -960 346748 480 346988 4 io_out[15]
port 141 nsew
rlabel metal2 s 58594 703520 58706 704960 6 io_out[16]
port 142 nsew
rlabel metal2 s 195766 703520 195878 704960 6 io_out[17]
port 143 nsew
rlabel metal2 s 23818 703520 23930 704960 6 io_out[18]
port 144 nsew
rlabel metal3 s 583520 266508 584960 266748 6 io_out[19]
port 145 nsew
rlabel metal3 s 583520 407268 584960 407508 6 io_out[1]
port 146 nsew
rlabel metal2 s 70186 703520 70298 704960 6 io_out[20]
port 147 nsew
rlabel metal2 s 271114 -960 271226 480 8 io_out[21]
port 148 nsew
rlabel metal3 s -960 184908 480 185148 4 io_out[22]
port 149 nsew
rlabel metal3 s 583520 354908 584960 355148 6 io_out[23]
port 150 nsew
rlabel metal3 s -960 685388 480 685628 4 io_out[24]
port 151 nsew
rlabel metal3 s -960 269908 480 270148 4 io_out[25]
port 152 nsew
rlabel metal2 s 221526 -960 221638 480 8 io_out[26]
port 153 nsew
rlabel metal2 s 179022 -960 179134 480 8 io_out[2]
port 154 nsew
rlabel metal2 s 276266 703520 276378 704960 6 io_out[3]
port 155 nsew
rlabel metal2 s 470754 703520 470866 704960 6 io_out[4]
port 156 nsew
rlabel metal3 s -960 483428 480 483668 4 io_out[5]
port 157 nsew
rlabel metal3 s 583520 165188 584960 165428 6 io_out[6]
port 158 nsew
rlabel metal3 s -960 653428 480 653668 4 io_out[7]
port 159 nsew
rlabel metal3 s 583520 120988 584960 121228 6 io_out[8]
port 160 nsew
rlabel metal3 s 583520 250188 584960 250428 6 io_out[9]
port 161 nsew
rlabel metal2 s 157770 703520 157882 704960 6 la_data_in[0]
port 162 nsew
rlabel metal3 s 583520 625548 584960 625788 6 la_data_in[100]
port 163 nsew
rlabel metal3 s 583520 214148 584960 214388 6 la_data_in[101]
port 164 nsew
rlabel metal2 s 387034 703520 387146 704960 6 la_data_in[102]
port 165 nsew
rlabel metal3 s 583520 20348 584960 20588 6 la_data_in[103]
port 166 nsew
rlabel metal3 s -960 370548 480 370788 4 la_data_in[104]
port 167 nsew
rlabel metal2 s 222814 703520 222926 704960 6 la_data_in[105]
port 168 nsew
rlabel metal2 s 134586 703520 134698 704960 6 la_data_in[106]
port 169 nsew
rlabel metal3 s -960 415428 480 415668 4 la_data_in[107]
port 170 nsew
rlabel metal3 s 583520 584748 584960 584988 6 la_data_in[108]
port 171 nsew
rlabel metal3 s -960 161108 480 161348 4 la_data_in[109]
port 172 nsew
rlabel metal3 s 583520 379388 584960 379628 6 la_data_in[10]
port 173 nsew
rlabel metal3 s -960 286228 480 286468 4 la_data_in[110]
port 174 nsew
rlabel metal3 s 583520 270588 584960 270828 6 la_data_in[111]
port 175 nsew
rlabel metal3 s -960 374628 480 374868 4 la_data_in[112]
port 176 nsew
rlabel metal3 s -960 673148 480 673388 4 la_data_in[113]
port 177 nsew
rlabel metal3 s -960 516068 480 516308 4 la_data_in[114]
port 178 nsew
rlabel metal2 s 325854 703520 325966 704960 6 la_data_in[115]
port 179 nsew
rlabel metal2 s 526782 -960 526894 480 8 la_data_in[116]
port 180 nsew
rlabel metal3 s -960 338588 480 338828 4 la_data_in[117]
port 181 nsew
rlabel metal3 s 583520 520828 584960 521068 6 la_data_in[118]
port 182 nsew
rlabel metal3 s 583520 210068 584960 210308 6 la_data_in[119]
port 183 nsew
rlabel metal2 s 96590 703520 96702 704960 6 la_data_in[11]
port 184 nsew
rlabel metal3 s -960 305948 480 306188 4 la_data_in[120]
port 185 nsew
rlabel metal2 s 160346 -960 160458 480 8 la_data_in[121]
port 186 nsew
rlabel metal2 s 137162 -960 137274 480 8 la_data_in[122]
port 187 nsew
rlabel metal3 s -960 426988 480 427228 4 la_data_in[123]
port 188 nsew
rlabel metal2 s 413438 703520 413550 704960 6 la_data_in[124]
port 189 nsew
rlabel metal2 s 484922 -960 485034 480 8 la_data_in[125]
port 190 nsew
rlabel metal3 s -960 419508 480 419748 4 la_data_in[126]
port 191 nsew
rlabel metal2 s 558982 703520 559094 704960 6 la_data_in[127]
port 192 nsew
rlabel metal3 s 583520 185588 584960 185828 6 la_data_in[12]
port 193 nsew
rlabel metal3 s 583520 339268 584960 339508 6 la_data_in[13]
port 194 nsew
rlabel metal3 s -960 539868 480 540108 4 la_data_in[14]
port 195 nsew
rlabel metal3 s -960 548028 480 548268 4 la_data_in[15]
port 196 nsew
rlabel metal3 s -960 67948 480 68188 4 la_data_in[16]
port 197 nsew
rlabel metal3 s -960 157028 480 157268 4 la_data_in[17]
port 198 nsew
rlabel metal3 s -960 451468 480 451708 4 la_data_in[18]
port 199 nsew
rlabel metal2 s 448214 703520 448326 704960 6 la_data_in[19]
port 200 nsew
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[1]
port 201 nsew
rlabel metal3 s -960 310028 480 310268 4 la_data_in[20]
port 202 nsew
rlabel metal2 s 27682 703520 27794 704960 6 la_data_in[21]
port 203 nsew
rlabel metal2 s 180954 703520 181066 704960 6 la_data_in[22]
port 204 nsew
rlabel metal3 s -960 439228 480 439468 4 la_data_in[23]
port 205 nsew
rlabel metal3 s 583520 423588 584960 423828 6 la_data_in[24]
port 206 nsew
rlabel metal2 s 432758 703520 432870 704960 6 la_data_in[25]
port 207 nsew
rlabel metal2 s 504242 -960 504354 480 8 la_data_in[26]
port 208 nsew
rlabel metal2 s 289790 -960 289902 480 8 la_data_in[27]
port 209 nsew
rlabel metal3 s -960 463708 480 463948 4 la_data_in[28]
port 210 nsew
rlabel metal3 s -960 342668 480 342908 4 la_data_in[29]
port 211 nsew
rlabel metal2 s 439198 -960 439310 480 8 la_data_in[2]
port 212 nsew
rlabel metal3 s -960 491588 480 491828 4 la_data_in[30]
port 213 nsew
rlabel metal3 s 583520 605148 584960 605388 6 la_data_in[31]
port 214 nsew
rlabel metal2 s 302670 703520 302782 704960 6 la_data_in[32]
port 215 nsew
rlabel metal3 s 583520 588828 584960 589068 6 la_data_in[33]
port 216 nsew
rlabel metal3 s -960 7428 480 7668 4 la_data_in[34]
port 217 nsew
rlabel metal3 s -960 664988 480 665228 4 la_data_in[35]
port 218 nsew
rlabel metal2 s 551254 703520 551366 704960 6 la_data_in[36]
port 219 nsew
rlabel metal2 s 543526 703520 543638 704960 6 la_data_in[37]
port 220 nsew
rlabel metal2 s 329718 703520 329830 704960 6 la_data_in[38]
port 221 nsew
rlabel metal2 s 148754 -960 148866 480 8 la_data_in[39]
port 222 nsew
rlabel metal3 s 583520 395708 584960 395948 6 la_data_in[3]
port 223 nsew
rlabel metal2 s 138450 703520 138562 704960 6 la_data_in[40]
port 224 nsew
rlabel metal3 s -960 620788 480 621028 4 la_data_in[41]
port 225 nsew
rlabel metal3 s -960 144788 480 145028 4 la_data_in[42]
port 226 nsew
rlabel metal3 s 583520 318868 584960 319108 6 la_data_in[43]
port 227 nsew
rlabel metal3 s -960 459628 480 459868 4 la_data_in[44]
port 228 nsew
rlabel metal2 s 81134 703520 81246 704960 6 la_data_in[45]
port 229 nsew
rlabel metal2 s 123638 703520 123750 704960 6 la_data_in[46]
port 230 nsew
rlabel metal3 s -960 580668 480 580908 4 la_data_in[47]
port 231 nsew
rlabel metal3 s 583520 419508 584960 419748 6 la_data_in[48]
port 232 nsew
rlabel metal3 s 583520 32588 584960 32828 6 la_data_in[49]
port 233 nsew
rlabel metal2 s 431470 -960 431582 480 8 la_data_in[4]
port 234 nsew
rlabel metal2 s 488786 -960 488898 480 8 la_data_in[50]
port 235 nsew
rlabel metal3 s 583520 500428 584960 500668 6 la_data_in[51]
port 236 nsew
rlabel metal3 s -960 552108 480 552348 4 la_data_in[52]
port 237 nsew
rlabel metal2 s 255658 -960 255770 480 8 la_data_in[53]
port 238 nsew
rlabel metal2 s 3210 -960 3322 480 8 la_data_in[54]
port 239 nsew
rlabel metal3 s 583520 322948 584960 323188 6 la_data_in[55]
port 240 nsew
rlabel metal3 s -960 507908 480 508148 4 la_data_in[56]
port 241 nsew
rlabel metal3 s 583520 411348 584960 411588 6 la_data_in[57]
port 242 nsew
rlabel metal2 s 394762 703520 394874 704960 6 la_data_in[58]
port 243 nsew
rlabel metal3 s -960 104668 480 104908 4 la_data_in[59]
port 244 nsew
rlabel metal3 s -960 612628 480 612868 4 la_data_in[5]
port 245 nsew
rlabel metal2 s 542238 -960 542350 480 8 la_data_in[60]
port 246 nsew
rlabel metal2 s 568642 -960 568754 480 8 la_data_in[61]
port 247 nsew
rlabel metal3 s 583520 48228 584960 48468 6 la_data_in[62]
port 248 nsew
rlabel metal3 s -960 188988 480 189228 4 la_data_in[63]
port 249 nsew
rlabel metal3 s 583520 173348 584960 173588 6 la_data_in[64]
port 250 nsew
rlabel metal3 s 583520 577268 584960 577508 6 la_data_in[65]
port 251 nsew
rlabel metal3 s 583520 331108 584960 331348 6 la_data_in[66]
port 252 nsew
rlabel metal2 s 79846 -960 79958 480 8 la_data_in[67]
port 253 nsew
rlabel metal3 s 583520 565028 584960 565268 6 la_data_in[68]
port 254 nsew
rlabel metal3 s 583520 677908 584960 678148 6 la_data_in[69]
port 255 nsew
rlabel metal3 s 583520 298468 584960 298708 6 la_data_in[6]
port 256 nsew
rlabel metal3 s -960 499748 480 499988 4 la_data_in[70]
port 257 nsew
rlabel metal3 s -960 165188 480 165428 4 la_data_in[71]
port 258 nsew
rlabel metal2 s 62458 703520 62570 704960 6 la_data_in[72]
port 259 nsew
rlabel metal3 s -960 100588 480 100828 4 la_data_in[73]
port 260 nsew
rlabel metal3 s 583520 327028 584960 327268 6 la_data_in[74]
port 261 nsew
rlabel metal2 s 127502 703520 127614 704960 6 la_data_in[75]
port 262 nsew
rlabel metal3 s 583520 149548 584960 149788 6 la_data_in[76]
port 263 nsew
rlabel metal2 s 165498 703520 165610 704960 6 la_data_in[77]
port 264 nsew
rlabel metal2 s 238270 703520 238382 704960 6 la_data_in[78]
port 265 nsew
rlabel metal3 s 583520 536468 584960 536708 6 la_data_in[79]
port 266 nsew
rlabel metal2 s 343242 -960 343354 480 8 la_data_in[7]
port 267 nsew
rlabel metal3 s -960 330428 480 330668 4 la_data_in[80]
port 268 nsew
rlabel metal2 s 505530 703520 505642 704960 6 la_data_in[81]
port 269 nsew
rlabel metal2 s 150042 703520 150154 704960 6 la_data_in[82]
port 270 nsew
rlabel metal3 s 583520 661588 584960 661828 6 la_data_in[83]
port 271 nsew
rlabel metal3 s -960 681308 480 681548 4 la_data_in[84]
port 272 nsew
rlabel metal3 s 583520 367148 584960 367388 6 la_data_in[85]
port 273 nsew
rlabel metal3 s 583520 448068 584960 448308 6 la_data_in[86]
port 274 nsew
rlabel metal2 s 95302 -960 95414 480 8 la_data_in[87]
port 275 nsew
rlabel metal3 s 583520 488188 584960 488428 6 la_data_in[88]
port 276 nsew
rlabel metal2 s 251794 -960 251906 480 8 la_data_in[89]
port 277 nsew
rlabel metal2 s 274978 -960 275090 480 8 la_data_in[8]
port 278 nsew
rlabel metal3 s -960 604468 480 604708 4 la_data_in[90]
port 279 nsew
rlabel metal3 s -960 532388 480 532628 4 la_data_in[91]
port 280 nsew
rlabel metal3 s 583520 12188 584960 12428 6 la_data_in[92]
port 281 nsew
rlabel metal3 s -960 197148 480 197388 4 la_data_in[93]
port 282 nsew
rlabel metal3 s 583520 314788 584960 315028 6 la_data_in[94]
port 283 nsew
rlabel metal3 s -960 96508 480 96748 4 la_data_in[95]
port 284 nsew
rlabel metal3 s -960 511988 480 512228 4 la_data_in[96]
port 285 nsew
rlabel metal3 s -960 568428 480 568668 4 la_data_in[97]
port 286 nsew
rlabel metal2 s 282706 -960 282818 480 8 la_data_in[98]
port 287 nsew
rlabel metal3 s 583520 573188 584960 573428 6 la_data_in[99]
port 288 nsew
rlabel metal2 s 119774 703520 119886 704960 6 la_data_in[9]
port 289 nsew
rlabel metal3 s -960 503828 480 504068 4 la_data_out[0]
port 290 nsew
rlabel metal2 s 253082 703520 253194 704960 6 la_data_out[100]
port 291 nsew
rlabel metal2 s 232474 -960 232586 480 8 la_data_out[101]
port 292 nsew
rlabel metal2 s 169362 703520 169474 704960 6 la_data_out[102]
port 293 nsew
rlabel metal3 s 583520 254268 584960 254508 6 la_data_out[103]
port 294 nsew
rlabel metal2 s 161634 703520 161746 704960 6 la_data_out[104]
port 295 nsew
rlabel metal3 s 583520 189668 584960 189908 6 la_data_out[105]
port 296 nsew
rlabel metal2 s 152618 -960 152730 480 8 la_data_out[106]
port 297 nsew
rlabel metal3 s 583520 387548 584960 387788 6 la_data_out[107]
port 298 nsew
rlabel metal3 s 583520 512668 584960 512908 6 la_data_out[108]
port 299 nsew
rlabel metal2 s 509394 703520 509506 704960 6 la_data_out[109]
port 300 nsew
rlabel metal3 s -960 386868 480 387108 4 la_data_out[10]
port 301 nsew
rlabel metal3 s -960 213468 480 213708 4 la_data_out[110]
port 302 nsew
rlabel metal3 s -960 282148 480 282388 4 la_data_out[111]
port 303 nsew
rlabel metal3 s -960 701708 480 701948 4 la_data_out[112]
port 304 nsew
rlabel metal2 s 202206 -960 202318 480 8 la_data_out[113]
port 305 nsew
rlabel metal2 s 570574 703520 570686 704960 6 la_data_out[114]
port 306 nsew
rlabel metal2 s 375442 703520 375554 704960 6 la_data_out[115]
port 307 nsew
rlabel metal2 s 408286 -960 408398 480 8 la_data_out[116]
port 308 nsew
rlabel metal3 s 583520 645268 584960 645508 6 la_data_out[117]
port 309 nsew
rlabel metal3 s 583520 391628 584960 391868 6 la_data_out[118]
port 310 nsew
rlabel metal3 s 583520 24428 584960 24668 6 la_data_out[119]
port 311 nsew
rlabel metal2 s 452078 703520 452190 704960 6 la_data_out[11]
port 312 nsew
rlabel metal2 s 18666 -960 18778 480 8 la_data_out[120]
port 313 nsew
rlabel metal2 s 184818 703520 184930 704960 6 la_data_out[121]
port 314 nsew
rlabel metal2 s 379306 703520 379418 704960 6 la_data_out[122]
port 315 nsew
rlabel metal3 s -960 229788 480 230028 4 la_data_out[123]
port 316 nsew
rlabel metal3 s 583520 137308 584960 137548 6 la_data_out[124]
port 317 nsew
rlabel metal3 s 583520 480028 584960 480268 6 la_data_out[125]
port 318 nsew
rlabel metal3 s -960 31908 480 32148 4 la_data_out[126]
port 319 nsew
rlabel metal3 s -960 354908 480 355148 4 la_data_out[127]
port 320 nsew
rlabel metal2 s 225390 -960 225502 480 8 la_data_out[12]
port 321 nsew
rlabel metal3 s 583520 40748 584960 40988 6 la_data_out[13]
port 322 nsew
rlabel metal3 s -960 362388 480 362628 4 la_data_out[14]
port 323 nsew
rlabel metal3 s -960 455548 480 455788 4 la_data_out[15]
port 324 nsew
rlabel metal2 s 341310 703520 341422 704960 6 la_data_out[16]
port 325 nsew
rlabel metal3 s 583520 431748 584960 431988 6 la_data_out[17]
port 326 nsew
rlabel metal2 s 110758 -960 110870 480 8 la_data_out[18]
port 327 nsew
rlabel metal2 s 188038 703520 188150 704960 6 la_data_out[19]
port 328 nsew
rlabel metal3 s 583520 93108 584960 93348 6 la_data_out[1]
port 329 nsew
rlabel metal3 s -960 27828 480 28068 4 la_data_out[20]
port 330 nsew
rlabel metal3 s 583520 225708 584960 225948 6 la_data_out[21]
port 331 nsew
rlabel metal3 s 583520 698308 584960 698548 6 la_data_out[22]
port 332 nsew
rlabel metal3 s 583520 229788 584960 230028 6 la_data_out[23]
port 333 nsew
rlabel metal3 s -960 689468 480 689708 4 la_data_out[24]
port 334 nsew
rlabel metal2 s 469466 -960 469578 480 8 la_data_out[25]
port 335 nsew
rlabel metal3 s 583520 467788 584960 468028 6 la_data_out[26]
port 336 nsew
rlabel metal3 s -960 92428 480 92668 4 la_data_out[27]
port 337 nsew
rlabel metal2 s 309110 -960 309222 480 8 la_data_out[28]
port 338 nsew
rlabel metal2 s 305246 -960 305358 480 8 la_data_out[29]
port 339 nsew
rlabel metal2 s 477194 -960 477306 480 8 la_data_out[2]
port 340 nsew
rlabel metal2 s 272402 703520 272514 704960 6 la_data_out[30]
port 341 nsew
rlabel metal3 s -960 237948 480 238188 4 la_data_out[31]
port 342 nsew
rlabel metal3 s -960 217548 480 217788 4 la_data_out[32]
port 343 nsew
rlabel metal3 s 583520 201908 584960 202148 6 la_data_out[33]
port 344 nsew
rlabel metal2 s 316838 -960 316950 480 8 la_data_out[34]
port 345 nsew
rlabel metal3 s -960 322268 480 322508 4 la_data_out[35]
port 346 nsew
rlabel metal2 s 528070 703520 528182 704960 6 la_data_out[36]
port 347 nsew
rlabel metal3 s 583520 8108 584960 8348 6 la_data_out[37]
port 348 nsew
rlabel metal3 s 583520 68628 584960 68868 6 la_data_out[38]
port 349 nsew
rlabel metal3 s 583520 129148 584960 129388 6 la_data_out[39]
port 350 nsew
rlabel metal3 s -960 80188 480 80428 4 la_data_out[3]
port 351 nsew
rlabel metal3 s 583520 346748 584960 346988 6 la_data_out[40]
port 352 nsew
rlabel metal2 s 371578 703520 371690 704960 6 la_data_out[41]
port 353 nsew
rlabel metal2 s 245354 703520 245466 704960 6 la_data_out[42]
port 354 nsew
rlabel metal3 s -960 693548 480 693788 4 la_data_out[43]
port 355 nsew
rlabel metal2 s 465602 -960 465714 480 8 la_data_out[44]
port 356 nsew
rlabel metal2 s 378018 -960 378130 480 8 la_data_out[45]
port 357 nsew
rlabel metal2 s 84998 703520 85110 704960 6 la_data_out[46]
port 358 nsew
rlabel metal3 s -960 628948 480 629188 4 la_data_out[47]
port 359 nsew
rlabel metal2 s 561558 -960 561670 480 8 la_data_out[48]
port 360 nsew
rlabel metal2 s 146178 703520 146290 704960 6 la_data_out[49]
port 361 nsew
rlabel metal2 s 486210 703520 486322 704960 6 la_data_out[4]
port 362 nsew
rlabel metal3 s -960 431068 480 431308 4 la_data_out[50]
port 363 nsew
rlabel metal2 s 370290 -960 370402 480 8 la_data_out[51]
port 364 nsew
rlabel metal3 s -960 84268 480 84508 4 la_data_out[52]
port 365 nsew
rlabel metal2 s 440486 703520 440598 704960 6 la_data_out[53]
port 366 nsew
rlabel metal2 s 397338 -960 397450 480 8 la_data_out[54]
port 367 nsew
rlabel metal3 s -960 201228 480 201468 4 la_data_out[55]
port 368 nsew
rlabel metal2 s 280130 703520 280242 704960 6 la_data_out[56]
port 369 nsew
rlabel metal2 s 47002 703520 47114 704960 6 la_data_out[57]
port 370 nsew
rlabel metal3 s 583520 125068 584960 125308 6 la_data_out[58]
port 371 nsew
rlabel metal3 s 583520 427668 584960 427908 6 la_data_out[59]
port 372 nsew
rlabel metal2 s 354834 -960 354946 480 8 la_data_out[5]
port 373 nsew
rlabel metal3 s -960 645268 480 645508 4 la_data_out[60]
port 374 nsew
rlabel metal3 s -960 411348 480 411588 4 la_data_out[61]
port 375 nsew
rlabel metal2 s 362562 -960 362674 480 8 la_data_out[62]
port 376 nsew
rlabel metal2 s 436622 703520 436734 704960 6 la_data_out[63]
port 377 nsew
rlabel metal3 s -960 273988 480 274228 4 la_data_out[64]
port 378 nsew
rlabel metal2 s 522918 -960 523030 480 8 la_data_out[65]
port 379 nsew
rlabel metal3 s 583520 -52 584960 188 6 la_data_out[66]
port 380 nsew
rlabel metal3 s -960 148868 480 149108 4 la_data_out[67]
port 381 nsew
rlabel metal3 s -960 63868 480 64108 4 la_data_out[68]
port 382 nsew
rlabel metal3 s 583520 181508 584960 181748 6 la_data_out[69]
port 383 nsew
rlabel metal2 s 320702 -960 320814 480 8 la_data_out[6]
port 384 nsew
rlabel metal2 s 473330 -960 473442 480 8 la_data_out[70]
port 385 nsew
rlabel metal3 s -960 48228 480 48468 4 la_data_out[71]
port 386 nsew
rlabel metal2 s 444350 703520 444462 704960 6 la_data_out[72]
port 387 nsew
rlabel metal2 s 358698 -960 358810 480 8 la_data_out[73]
port 388 nsew
rlabel metal2 s 5142 703520 5254 704960 6 la_data_out[74]
port 389 nsew
rlabel metal2 s 400558 -960 400670 480 8 la_data_out[75]
port 390 nsew
rlabel metal3 s -960 669068 480 669308 4 la_data_out[76]
port 391 nsew
rlabel metal3 s 583520 475948 584960 476188 6 la_data_out[77]
port 392 nsew
rlabel metal2 s 332294 -960 332406 480 8 la_data_out[78]
port 393 nsew
rlabel metal3 s 583520 153628 584960 153868 6 la_data_out[79]
port 394 nsew
rlabel metal3 s 583520 44148 584960 44388 6 la_data_out[7]
port 395 nsew
rlabel metal3 s 583520 233868 584960 234108 6 la_data_out[80]
port 396 nsew
rlabel metal3 s -960 572508 480 572748 4 la_data_out[81]
port 397 nsew
rlabel metal2 s 247930 -960 248042 480 8 la_data_out[82]
port 398 nsew
rlabel metal3 s -960 560268 480 560508 4 la_data_out[83]
port 399 nsew
rlabel metal2 s 461738 -960 461850 480 8 la_data_out[84]
port 400 nsew
rlabel metal2 s 517122 703520 517234 704960 6 la_data_out[85]
port 401 nsew
rlabel metal2 s 115910 703520 116022 704960 6 la_data_out[86]
port 402 nsew
rlabel metal2 s 578302 703520 578414 704960 6 la_data_out[87]
port 403 nsew
rlabel metal3 s -960 112828 480 113068 4 la_data_out[88]
port 404 nsew
rlabel metal3 s 583520 76788 584960 77028 6 la_data_out[89]
port 405 nsew
rlabel metal3 s 583520 439908 584960 440148 6 la_data_out[8]
port 406 nsew
rlabel metal2 s 226678 703520 226790 704960 6 la_data_out[90]
port 407 nsew
rlabel metal2 s 423742 -960 423854 480 8 la_data_out[91]
port 408 nsew
rlabel metal2 s 171294 -960 171406 480 8 la_data_out[92]
port 409 nsew
rlabel metal2 s 417302 703520 417414 704960 6 la_data_out[93]
port 410 nsew
rlabel metal2 s 496514 -960 496626 480 8 la_data_out[94]
port 411 nsew
rlabel metal3 s -960 278068 480 278308 4 la_data_out[95]
port 412 nsew
rlabel metal2 s 9006 703520 9118 704960 6 la_data_out[96]
port 413 nsew
rlabel metal2 s 190614 -960 190726 480 8 la_data_out[97]
port 414 nsew
rlabel metal2 s 555118 703520 555230 704960 6 la_data_out[98]
port 415 nsew
rlabel metal2 s 511326 -960 511438 480 8 la_data_out[99]
port 416 nsew
rlabel metal3 s 583520 286228 584960 286468 6 la_data_out[9]
port 417 nsew
rlabel metal2 s 425030 703520 425142 704960 6 la_oenb[0]
port 418 nsew
rlabel metal3 s -960 209388 480 209628 4 la_oenb[100]
port 419 nsew
rlabel metal3 s -960 480028 480 480268 4 la_oenb[101]
port 420 nsew
rlabel metal2 s 297518 -960 297630 480 8 la_oenb[102]
port 421 nsew
rlabel metal2 s 350970 -960 351082 480 8 la_oenb[103]
port 422 nsew
rlabel metal2 s 43138 703520 43250 704960 6 la_oenb[104]
port 423 nsew
rlabel metal3 s 583520 161788 584960 162028 6 la_oenb[105]
port 424 nsew
rlabel metal2 s 421166 703520 421278 704960 6 la_oenb[106]
port 425 nsew
rlabel metal2 s 168074 -960 168186 480 8 la_oenb[107]
port 426 nsew
rlabel metal3 s 583520 471868 584960 472108 6 la_oenb[108]
port 427 nsew
rlabel metal2 s 177090 703520 177202 704960 6 la_oenb[109]
port 428 nsew
rlabel metal2 s 513258 703520 513370 704960 6 la_oenb[10]
port 429 nsew
rlabel metal2 s 142314 703520 142426 704960 6 la_oenb[110]
port 430 nsew
rlabel metal2 s 35410 703520 35522 704960 6 la_oenb[111]
port 431 nsew
rlabel metal3 s -960 120308 480 120548 4 la_oenb[112]
port 432 nsew
rlabel metal2 s 263386 -960 263498 480 8 la_oenb[113]
port 433 nsew
rlabel metal3 s 583520 596988 584960 597228 6 la_oenb[114]
port 434 nsew
rlabel metal2 s 481058 -960 481170 480 8 la_oenb[115]
port 435 nsew
rlabel metal3 s 583520 435828 584960 436068 6 la_oenb[116]
port 436 nsew
rlabel metal2 s 125570 -960 125682 480 8 la_oenb[117]
port 437 nsew
rlabel metal2 s 260810 703520 260922 704960 6 la_oenb[118]
port 438 nsew
rlabel metal3 s -960 44148 480 44388 4 la_oenb[119]
port 439 nsew
rlabel metal2 s 340022 -960 340134 480 8 la_oenb[11]
port 440 nsew
rlabel metal2 s 562846 703520 562958 704960 6 la_oenb[120]
port 441 nsew
rlabel metal3 s -960 378708 480 378948 4 la_oenb[121]
port 442 nsew
rlabel metal3 s 583520 112828 584960 113068 6 la_oenb[122]
port 443 nsew
rlabel metal2 s 12870 703520 12982 704960 6 la_oenb[123]
port 444 nsew
rlabel metal2 s 50866 703520 50978 704960 6 la_oenb[124]
port 445 nsew
rlabel metal2 s 236338 -960 236450 480 8 la_oenb[125]
port 446 nsew
rlabel metal2 s 287858 703520 287970 704960 6 la_oenb[126]
port 447 nsew
rlabel metal3 s 583520 637788 584960 638028 6 la_oenb[127]
port 448 nsew
rlabel metal3 s 583520 302548 584960 302788 6 la_oenb[12]
port 449 nsew
rlabel metal3 s -960 318188 480 318428 4 la_oenb[13]
port 450 nsew
rlabel metal3 s -960 193068 480 193308 4 la_oenb[14]
port 451 nsew
rlabel metal3 s 583520 246108 584960 246348 6 la_oenb[15]
port 452 nsew
rlabel metal3 s -960 40068 480 40308 4 la_oenb[16]
port 453 nsew
rlabel metal2 s 283994 703520 284106 704960 6 la_oenb[17]
port 454 nsew
rlabel metal3 s -960 152948 480 153188 4 la_oenb[18]
port 455 nsew
rlabel metal3 s -960 72028 480 72268 4 la_oenb[19]
port 456 nsew
rlabel metal2 s 186750 -960 186862 480 8 la_oenb[1]
port 457 nsew
rlabel metal3 s 583520 193748 584960 193988 6 la_oenb[20]
port 458 nsew
rlabel metal2 s 41850 -960 41962 480 8 la_oenb[21]
port 459 nsew
rlabel metal2 s 194478 -960 194590 480 8 la_oenb[22]
port 460 nsew
rlabel metal3 s 583520 177428 584960 177668 6 la_oenb[23]
port 461 nsew
rlabel metal2 s 582166 703520 582278 704960 6 la_oenb[24]
port 462 nsew
rlabel metal3 s 583520 358988 584960 359228 6 la_oenb[25]
port 463 nsew
rlabel metal2 s 68254 -960 68366 480 8 la_oenb[26]
port 464 nsew
rlabel metal3 s 583520 306628 584960 306868 6 la_oenb[27]
port 465 nsew
rlabel metal3 s -960 15588 480 15828 4 la_oenb[28]
port 466 nsew
rlabel metal2 s 459806 703520 459918 704960 6 la_oenb[29]
port 467 nsew
rlabel metal2 s 419878 -960 419990 480 8 la_oenb[2]
port 468 nsew
rlabel metal3 s 583520 443988 584960 444228 6 la_oenb[30]
port 469 nsew
rlabel metal2 s 539662 703520 539774 704960 6 la_oenb[31]
port 470 nsew
rlabel metal3 s -960 23748 480 23988 4 la_oenb[32]
port 471 nsew
rlabel metal2 s 306534 703520 306646 704960 6 la_oenb[33]
port 472 nsew
rlabel metal2 s 547390 703520 547502 704960 6 la_oenb[34]
port 473 nsew
rlabel metal2 s 77270 703520 77382 704960 6 la_oenb[35]
port 474 nsew
rlabel metal3 s -960 301868 480 302108 4 la_oenb[36]
port 475 nsew
rlabel metal3 s 583520 116908 584960 117148 6 la_oenb[37]
port 476 nsew
rlabel metal3 s -960 290308 480 290548 4 la_oenb[38]
port 477 nsew
rlabel metal3 s 583520 463708 584960 463948 6 la_oenb[39]
port 478 nsew
rlabel metal2 s 215086 703520 215198 704960 6 la_oenb[3]
port 479 nsew
rlabel metal2 s 500378 -960 500490 480 8 la_oenb[40]
port 480 nsew
rlabel metal3 s 583520 617388 584960 617628 6 la_oenb[41]
port 481 nsew
rlabel metal3 s 583520 532388 584960 532628 6 la_oenb[42]
port 482 nsew
rlabel metal2 s 490074 703520 490186 704960 6 la_oenb[43]
port 483 nsew
rlabel metal3 s 583520 681988 584960 682228 6 la_oenb[44]
port 484 nsew
rlabel metal3 s 583520 16268 584960 16508 6 la_oenb[45]
port 485 nsew
rlabel metal3 s -960 11508 480 11748 4 la_oenb[46]
port 486 nsew
rlabel metal2 s 576370 -960 576482 480 8 la_oenb[47]
port 487 nsew
rlabel metal3 s 583520 108748 584960 108988 6 la_oenb[48]
port 488 nsew
rlabel metal2 s 117842 -960 117954 480 8 la_oenb[49]
port 489 nsew
rlabel metal2 s 175158 -960 175270 480 8 la_oenb[4]
port 490 nsew
rlabel metal3 s 583520 36668 584960 36908 6 la_oenb[50]
port 491 nsew
rlabel metal3 s 583520 274668 584960 274908 6 la_oenb[51]
port 492 nsew
rlabel metal3 s 583520 621468 584960 621708 6 la_oenb[52]
port 493 nsew
rlabel metal2 s 234406 703520 234518 704960 6 la_oenb[53]
port 494 nsew
rlabel metal2 s 203494 703520 203606 704960 6 la_oenb[54]
port 495 nsew
rlabel metal2 s 104318 703520 104430 704960 6 la_oenb[55]
port 496 nsew
rlabel metal2 s 217662 -960 217774 480 8 la_oenb[56]
port 497 nsew
rlabel metal3 s 583520 690148 584960 690388 6 la_oenb[57]
port 498 nsew
rlabel metal3 s -960 180828 480 181068 4 la_oenb[58]
port 499 nsew
rlabel metal2 s 66322 703520 66434 704960 6 la_oenb[59]
port 500 nsew
rlabel metal3 s -960 52308 480 52548 4 la_oenb[5]
port 501 nsew
rlabel metal3 s 583520 609228 584960 609468 6 la_oenb[60]
port 502 nsew
rlabel metal2 s 356122 703520 356234 704960 6 la_oenb[61]
port 503 nsew
rlabel metal2 s 314262 703520 314374 704960 6 la_oenb[62]
port 504 nsew
rlabel metal2 s 428894 703520 429006 704960 6 la_oenb[63]
port 505 nsew
rlabel metal2 s 463670 703520 463782 704960 6 la_oenb[64]
port 506 nsew
rlabel metal2 s 467534 703520 467646 704960 6 la_oenb[65]
port 507 nsew
rlabel metal3 s -960 241348 480 241588 4 la_oenb[66]
port 508 nsew
rlabel metal2 s 249218 703520 249330 704960 6 la_oenb[67]
port 509 nsew
rlabel metal3 s -960 225708 480 225948 4 la_oenb[68]
port 510 nsew
rlabel metal2 s 7074 -960 7186 480 8 la_oenb[69]
port 511 nsew
rlabel metal2 s 572506 -960 572618 480 8 la_oenb[6]
port 512 nsew
rlabel metal3 s -960 253588 480 253828 4 la_oenb[70]
port 513 nsew
rlabel metal3 s 583520 197828 584960 198068 6 la_oenb[71]
port 514 nsew
rlabel metal3 s -960 443308 480 443548 4 la_oenb[72]
port 515 nsew
rlabel metal3 s 583520 262428 584960 262668 6 la_oenb[73]
port 516 nsew
rlabel metal3 s -960 584748 480 584988 4 la_oenb[74]
port 517 nsew
rlabel metal2 s 30258 -960 30370 480 8 la_oenb[75]
port 518 nsew
rlabel metal3 s -960 261748 480 261988 4 la_oenb[76]
port 519 nsew
rlabel metal3 s -960 173348 480 173588 4 la_oenb[77]
port 520 nsew
rlabel metal2 s 242134 703520 242246 704960 6 la_oenb[78]
port 521 nsew
rlabel metal3 s 583520 4028 584960 4268 6 la_oenb[79]
port 522 nsew
rlabel metal2 s 278842 -960 278954 480 8 la_oenb[7]
port 523 nsew
rlabel metal3 s -960 495668 480 495908 4 la_oenb[80]
port 524 nsew
rlabel metal3 s 583520 528308 584960 528548 6 la_oenb[81]
port 525 nsew
rlabel metal3 s 583520 669748 584960 669988 6 la_oenb[82]
port 526 nsew
rlabel metal2 s 565422 -960 565534 480 8 la_oenb[83]
port 527 nsew
rlabel metal3 s -960 588828 480 589068 4 la_oenb[84]
port 528 nsew
rlabel metal3 s 583520 141388 584960 141628 6 la_oenb[85]
port 529 nsew
rlabel metal3 s 583520 633708 584960 633948 6 la_oenb[86]
port 530 nsew
rlabel metal2 s 153906 703520 154018 704960 6 la_oenb[87]
port 531 nsew
rlabel metal3 s 583520 540548 584960 540788 6 la_oenb[88]
port 532 nsew
rlabel metal2 s 549966 -960 550078 480 8 la_oenb[89]
port 533 nsew
rlabel metal2 s 310398 703520 310510 704960 6 la_oenb[8]
port 534 nsew
rlabel metal3 s 583520 218228 584960 218468 6 la_oenb[90]
port 535 nsew
rlabel metal2 s 108182 703520 108294 704960 6 la_oenb[91]
port 536 nsew
rlabel metal3 s 583520 84948 584960 85188 6 la_oenb[92]
port 537 nsew
rlabel metal3 s -960 422908 480 423148 4 la_oenb[93]
port 538 nsew
rlabel metal2 s 91438 -960 91550 480 8 la_oenb[94]
port 539 nsew
rlabel metal3 s 583520 516748 584960 516988 6 la_oenb[95]
port 540 nsew
rlabel metal2 s 404422 -960 404534 480 8 la_oenb[96]
port 541 nsew
rlabel metal3 s -960 221628 480 221868 4 la_oenb[97]
port 542 nsew
rlabel metal2 s 182886 -960 182998 480 8 la_oenb[98]
port 543 nsew
rlabel metal3 s -960 294388 480 294628 4 la_oenb[99]
port 544 nsew
rlabel metal3 s -960 616708 480 616948 4 la_oenb[9]
port 545 nsew
rlabel metal2 s 318126 703520 318238 704960 6 user_clock2
port 546 nsew
rlabel metal3 s 583520 702388 584960 702628 6 user_irq[0]
port 547 nsew
rlabel metal3 s -960 596988 480 597228 4 user_irq[1]
port 548 nsew
rlabel metal3 s -960 660908 480 661148 4 user_irq[2]
port 549 nsew
rlabel metal5 s -8726 686866 592650 687486 6 vccd1
port 550 nsew
rlabel metal5 s -8726 650866 592650 651486 6 vccd1
port 550 nsew
rlabel metal5 s -8726 614866 592650 615486 6 vccd1
port 550 nsew
rlabel metal5 s -8726 578866 592650 579486 6 vccd1
port 550 nsew
rlabel metal5 s -8726 542866 592650 543486 6 vccd1
port 550 nsew
rlabel metal5 s -8726 506866 592650 507486 6 vccd1
port 550 nsew
rlabel metal5 s -8726 470866 592650 471486 6 vccd1
port 550 nsew
rlabel metal5 s -8726 434866 592650 435486 6 vccd1
port 550 nsew
rlabel metal5 s -8726 398866 592650 399486 6 vccd1
port 550 nsew
rlabel metal5 s -8726 362866 592650 363486 6 vccd1
port 550 nsew
rlabel metal5 s -8726 326866 592650 327486 6 vccd1
port 550 nsew
rlabel metal5 s -8726 290866 592650 291486 6 vccd1
port 550 nsew
rlabel metal5 s -8726 254866 592650 255486 6 vccd1
port 550 nsew
rlabel metal5 s -8726 218866 592650 219486 6 vccd1
port 550 nsew
rlabel metal5 s -8726 182866 592650 183486 6 vccd1
port 550 nsew
rlabel metal5 s -8726 146866 592650 147486 6 vccd1
port 550 nsew
rlabel metal5 s -8726 110866 592650 111486 6 vccd1
port 550 nsew
rlabel metal5 s -8726 74866 592650 75486 6 vccd1
port 550 nsew
rlabel metal5 s -8726 38866 592650 39486 6 vccd1
port 550 nsew
rlabel metal5 s -8726 2866 592650 3486 6 vccd1
port 550 nsew
rlabel metal4 s 577794 -7654 578414 711590 6 vccd1
port 550 nsew
rlabel metal4 s 541794 -7654 542414 711590 6 vccd1
port 550 nsew
rlabel metal4 s 505794 -7654 506414 711590 6 vccd1
port 550 nsew
rlabel metal4 s 469794 -7654 470414 711590 6 vccd1
port 550 nsew
rlabel metal4 s 433794 -7654 434414 711590 6 vccd1
port 550 nsew
rlabel metal4 s 397794 -7654 398414 711590 6 vccd1
port 550 nsew
rlabel metal4 s 361794 -7654 362414 711590 6 vccd1
port 550 nsew
rlabel metal4 s 325794 -7654 326414 711590 6 vccd1
port 550 nsew
rlabel metal4 s 289794 -7654 290414 711590 6 vccd1
port 550 nsew
rlabel metal4 s 253794 -7654 254414 711590 6 vccd1
port 550 nsew
rlabel metal4 s 217794 -7654 218414 711590 6 vccd1
port 550 nsew
rlabel metal4 s 181794 -7654 182414 711590 6 vccd1
port 550 nsew
rlabel metal4 s 145794 -7654 146414 711590 6 vccd1
port 550 nsew
rlabel metal4 s 109794 -7654 110414 711590 6 vccd1
port 550 nsew
rlabel metal4 s 73794 -7654 74414 711590 6 vccd1
port 550 nsew
rlabel metal4 s 37794 -7654 38414 711590 6 vccd1
port 550 nsew
rlabel metal4 s 1794 -7654 2414 711590 6 vccd1
port 550 nsew
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 550 nsew
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 550 nsew
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 550 nsew
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 550 nsew
rlabel metal5 s -8726 694306 592650 694926 6 vccd2
port 551 nsew
rlabel metal5 s -8726 658306 592650 658926 6 vccd2
port 551 nsew
rlabel metal5 s -8726 622306 592650 622926 6 vccd2
port 551 nsew
rlabel metal5 s -8726 586306 592650 586926 6 vccd2
port 551 nsew
rlabel metal5 s -8726 550306 592650 550926 6 vccd2
port 551 nsew
rlabel metal5 s -8726 514306 592650 514926 6 vccd2
port 551 nsew
rlabel metal5 s -8726 478306 592650 478926 6 vccd2
port 551 nsew
rlabel metal5 s -8726 442306 592650 442926 6 vccd2
port 551 nsew
rlabel metal5 s -8726 406306 592650 406926 6 vccd2
port 551 nsew
rlabel metal5 s -8726 370306 592650 370926 6 vccd2
port 551 nsew
rlabel metal5 s -8726 334306 592650 334926 6 vccd2
port 551 nsew
rlabel metal5 s -8726 298306 592650 298926 6 vccd2
port 551 nsew
rlabel metal5 s -8726 262306 592650 262926 6 vccd2
port 551 nsew
rlabel metal5 s -8726 226306 592650 226926 6 vccd2
port 551 nsew
rlabel metal5 s -8726 190306 592650 190926 6 vccd2
port 551 nsew
rlabel metal5 s -8726 154306 592650 154926 6 vccd2
port 551 nsew
rlabel metal5 s -8726 118306 592650 118926 6 vccd2
port 551 nsew
rlabel metal5 s -8726 82306 592650 82926 6 vccd2
port 551 nsew
rlabel metal5 s -8726 46306 592650 46926 6 vccd2
port 551 nsew
rlabel metal5 s -8726 10306 592650 10926 6 vccd2
port 551 nsew
rlabel metal4 s 549234 -7654 549854 711590 6 vccd2
port 551 nsew
rlabel metal4 s 513234 -7654 513854 711590 6 vccd2
port 551 nsew
rlabel metal4 s 477234 -7654 477854 711590 6 vccd2
port 551 nsew
rlabel metal4 s 441234 -7654 441854 711590 6 vccd2
port 551 nsew
rlabel metal4 s 405234 -7654 405854 711590 6 vccd2
port 551 nsew
rlabel metal4 s 369234 -7654 369854 711590 6 vccd2
port 551 nsew
rlabel metal4 s 333234 -7654 333854 711590 6 vccd2
port 551 nsew
rlabel metal4 s 297234 -7654 297854 711590 6 vccd2
port 551 nsew
rlabel metal4 s 261234 -7654 261854 711590 6 vccd2
port 551 nsew
rlabel metal4 s 225234 -7654 225854 711590 6 vccd2
port 551 nsew
rlabel metal4 s 189234 -7654 189854 711590 6 vccd2
port 551 nsew
rlabel metal4 s 153234 -7654 153854 711590 6 vccd2
port 551 nsew
rlabel metal4 s 117234 -7654 117854 711590 6 vccd2
port 551 nsew
rlabel metal4 s 81234 -7654 81854 711590 6 vccd2
port 551 nsew
rlabel metal4 s 45234 -7654 45854 711590 6 vccd2
port 551 nsew
rlabel metal4 s 9234 -7654 9854 711590 6 vccd2
port 551 nsew
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 551 nsew
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 551 nsew
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 551 nsew
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 551 nsew
rlabel metal5 s -8726 665746 592650 666366 6 vdda1
port 552 nsew
rlabel metal5 s -8726 629746 592650 630366 6 vdda1
port 552 nsew
rlabel metal5 s -8726 593746 592650 594366 6 vdda1
port 552 nsew
rlabel metal5 s -8726 557746 592650 558366 6 vdda1
port 552 nsew
rlabel metal5 s -8726 521746 592650 522366 6 vdda1
port 552 nsew
rlabel metal5 s -8726 485746 592650 486366 6 vdda1
port 552 nsew
rlabel metal5 s -8726 449746 592650 450366 6 vdda1
port 552 nsew
rlabel metal5 s -8726 413746 592650 414366 6 vdda1
port 552 nsew
rlabel metal5 s -8726 377746 592650 378366 6 vdda1
port 552 nsew
rlabel metal5 s -8726 341746 592650 342366 6 vdda1
port 552 nsew
rlabel metal5 s -8726 305746 592650 306366 6 vdda1
port 552 nsew
rlabel metal5 s -8726 269746 592650 270366 6 vdda1
port 552 nsew
rlabel metal5 s -8726 233746 592650 234366 6 vdda1
port 552 nsew
rlabel metal5 s -8726 197746 592650 198366 6 vdda1
port 552 nsew
rlabel metal5 s -8726 161746 592650 162366 6 vdda1
port 552 nsew
rlabel metal5 s -8726 125746 592650 126366 6 vdda1
port 552 nsew
rlabel metal5 s -8726 89746 592650 90366 6 vdda1
port 552 nsew
rlabel metal5 s -8726 53746 592650 54366 6 vdda1
port 552 nsew
rlabel metal5 s -8726 17746 592650 18366 6 vdda1
port 552 nsew
rlabel metal4 s 556674 -7654 557294 711590 6 vdda1
port 552 nsew
rlabel metal4 s 520674 -7654 521294 711590 6 vdda1
port 552 nsew
rlabel metal4 s 484674 -7654 485294 711590 6 vdda1
port 552 nsew
rlabel metal4 s 448674 -7654 449294 711590 6 vdda1
port 552 nsew
rlabel metal4 s 412674 -7654 413294 711590 6 vdda1
port 552 nsew
rlabel metal4 s 376674 -7654 377294 711590 6 vdda1
port 552 nsew
rlabel metal4 s 340674 -7654 341294 711590 6 vdda1
port 552 nsew
rlabel metal4 s 304674 -7654 305294 711590 6 vdda1
port 552 nsew
rlabel metal4 s 268674 -7654 269294 711590 6 vdda1
port 552 nsew
rlabel metal4 s 232674 -7654 233294 711590 6 vdda1
port 552 nsew
rlabel metal4 s 196674 -7654 197294 711590 6 vdda1
port 552 nsew
rlabel metal4 s 160674 -7654 161294 711590 6 vdda1
port 552 nsew
rlabel metal4 s 124674 -7654 125294 711590 6 vdda1
port 552 nsew
rlabel metal4 s 88674 -7654 89294 711590 6 vdda1
port 552 nsew
rlabel metal4 s 52674 -7654 53294 711590 6 vdda1
port 552 nsew
rlabel metal4 s 16674 -7654 17294 711590 6 vdda1
port 552 nsew
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 552 nsew
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 552 nsew
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 552 nsew
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 552 nsew
rlabel metal5 s -8726 673186 592650 673806 6 vdda2
port 553 nsew
rlabel metal5 s -8726 637186 592650 637806 6 vdda2
port 553 nsew
rlabel metal5 s -8726 601186 592650 601806 6 vdda2
port 553 nsew
rlabel metal5 s -8726 565186 592650 565806 6 vdda2
port 553 nsew
rlabel metal5 s -8726 529186 592650 529806 6 vdda2
port 553 nsew
rlabel metal5 s -8726 493186 592650 493806 6 vdda2
port 553 nsew
rlabel metal5 s -8726 457186 592650 457806 6 vdda2
port 553 nsew
rlabel metal5 s -8726 421186 592650 421806 6 vdda2
port 553 nsew
rlabel metal5 s -8726 385186 592650 385806 6 vdda2
port 553 nsew
rlabel metal5 s -8726 349186 592650 349806 6 vdda2
port 553 nsew
rlabel metal5 s -8726 313186 592650 313806 6 vdda2
port 553 nsew
rlabel metal5 s -8726 277186 592650 277806 6 vdda2
port 553 nsew
rlabel metal5 s -8726 241186 592650 241806 6 vdda2
port 553 nsew
rlabel metal5 s -8726 205186 592650 205806 6 vdda2
port 553 nsew
rlabel metal5 s -8726 169186 592650 169806 6 vdda2
port 553 nsew
rlabel metal5 s -8726 133186 592650 133806 6 vdda2
port 553 nsew
rlabel metal5 s -8726 97186 592650 97806 6 vdda2
port 553 nsew
rlabel metal5 s -8726 61186 592650 61806 6 vdda2
port 553 nsew
rlabel metal5 s -8726 25186 592650 25806 6 vdda2
port 553 nsew
rlabel metal4 s 564114 -7654 564734 711590 6 vdda2
port 553 nsew
rlabel metal4 s 528114 -7654 528734 711590 6 vdda2
port 553 nsew
rlabel metal4 s 492114 -7654 492734 711590 6 vdda2
port 553 nsew
rlabel metal4 s 456114 -7654 456734 711590 6 vdda2
port 553 nsew
rlabel metal4 s 420114 -7654 420734 711590 6 vdda2
port 553 nsew
rlabel metal4 s 384114 -7654 384734 711590 6 vdda2
port 553 nsew
rlabel metal4 s 348114 -7654 348734 711590 6 vdda2
port 553 nsew
rlabel metal4 s 312114 -7654 312734 711590 6 vdda2
port 553 nsew
rlabel metal4 s 276114 -7654 276734 711590 6 vdda2
port 553 nsew
rlabel metal4 s 240114 -7654 240734 711590 6 vdda2
port 553 nsew
rlabel metal4 s 204114 -7654 204734 711590 6 vdda2
port 553 nsew
rlabel metal4 s 168114 -7654 168734 711590 6 vdda2
port 553 nsew
rlabel metal4 s 132114 -7654 132734 711590 6 vdda2
port 553 nsew
rlabel metal4 s 96114 -7654 96734 711590 6 vdda2
port 553 nsew
rlabel metal4 s 60114 -7654 60734 711590 6 vdda2
port 553 nsew
rlabel metal4 s 24114 -7654 24734 711590 6 vdda2
port 553 nsew
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 553 nsew
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 553 nsew
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 553 nsew
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 553 nsew
rlabel metal5 s -8726 669466 592650 670086 6 vssa1
port 554 nsew
rlabel metal5 s -8726 633466 592650 634086 6 vssa1
port 554 nsew
rlabel metal5 s -8726 597466 592650 598086 6 vssa1
port 554 nsew
rlabel metal5 s -8726 561466 592650 562086 6 vssa1
port 554 nsew
rlabel metal5 s -8726 525466 592650 526086 6 vssa1
port 554 nsew
rlabel metal5 s -8726 489466 592650 490086 6 vssa1
port 554 nsew
rlabel metal5 s -8726 453466 592650 454086 6 vssa1
port 554 nsew
rlabel metal5 s -8726 417466 592650 418086 6 vssa1
port 554 nsew
rlabel metal5 s -8726 381466 592650 382086 6 vssa1
port 554 nsew
rlabel metal5 s -8726 345466 592650 346086 6 vssa1
port 554 nsew
rlabel metal5 s -8726 309466 592650 310086 6 vssa1
port 554 nsew
rlabel metal5 s -8726 273466 592650 274086 6 vssa1
port 554 nsew
rlabel metal5 s -8726 237466 592650 238086 6 vssa1
port 554 nsew
rlabel metal5 s -8726 201466 592650 202086 6 vssa1
port 554 nsew
rlabel metal5 s -8726 165466 592650 166086 6 vssa1
port 554 nsew
rlabel metal5 s -8726 129466 592650 130086 6 vssa1
port 554 nsew
rlabel metal5 s -8726 93466 592650 94086 6 vssa1
port 554 nsew
rlabel metal5 s -8726 57466 592650 58086 6 vssa1
port 554 nsew
rlabel metal5 s -8726 21466 592650 22086 6 vssa1
port 554 nsew
rlabel metal4 s 560394 -7654 561014 711590 6 vssa1
port 554 nsew
rlabel metal4 s 524394 -7654 525014 711590 6 vssa1
port 554 nsew
rlabel metal4 s 488394 -7654 489014 711590 6 vssa1
port 554 nsew
rlabel metal4 s 452394 -7654 453014 711590 6 vssa1
port 554 nsew
rlabel metal4 s 416394 -7654 417014 711590 6 vssa1
port 554 nsew
rlabel metal4 s 380394 -7654 381014 711590 6 vssa1
port 554 nsew
rlabel metal4 s 344394 -7654 345014 711590 6 vssa1
port 554 nsew
rlabel metal4 s 308394 -7654 309014 711590 6 vssa1
port 554 nsew
rlabel metal4 s 272394 -7654 273014 711590 6 vssa1
port 554 nsew
rlabel metal4 s 236394 -7654 237014 711590 6 vssa1
port 554 nsew
rlabel metal4 s 200394 -7654 201014 711590 6 vssa1
port 554 nsew
rlabel metal4 s 164394 -7654 165014 711590 6 vssa1
port 554 nsew
rlabel metal4 s 128394 -7654 129014 711590 6 vssa1
port 554 nsew
rlabel metal4 s 92394 -7654 93014 711590 6 vssa1
port 554 nsew
rlabel metal4 s 56394 -7654 57014 711590 6 vssa1
port 554 nsew
rlabel metal4 s 20394 -7654 21014 711590 6 vssa1
port 554 nsew
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 554 nsew
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 554 nsew
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 554 nsew
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 554 nsew
rlabel metal5 s -8726 676906 592650 677526 6 vssa2
port 555 nsew
rlabel metal5 s -8726 640906 592650 641526 6 vssa2
port 555 nsew
rlabel metal5 s -8726 604906 592650 605526 6 vssa2
port 555 nsew
rlabel metal5 s -8726 568906 592650 569526 6 vssa2
port 555 nsew
rlabel metal5 s -8726 532906 592650 533526 6 vssa2
port 555 nsew
rlabel metal5 s -8726 496906 592650 497526 6 vssa2
port 555 nsew
rlabel metal5 s -8726 460906 592650 461526 6 vssa2
port 555 nsew
rlabel metal5 s -8726 424906 592650 425526 6 vssa2
port 555 nsew
rlabel metal5 s -8726 388906 592650 389526 6 vssa2
port 555 nsew
rlabel metal5 s -8726 352906 592650 353526 6 vssa2
port 555 nsew
rlabel metal5 s -8726 316906 592650 317526 6 vssa2
port 555 nsew
rlabel metal5 s -8726 280906 592650 281526 6 vssa2
port 555 nsew
rlabel metal5 s -8726 244906 592650 245526 6 vssa2
port 555 nsew
rlabel metal5 s -8726 208906 592650 209526 6 vssa2
port 555 nsew
rlabel metal5 s -8726 172906 592650 173526 6 vssa2
port 555 nsew
rlabel metal5 s -8726 136906 592650 137526 6 vssa2
port 555 nsew
rlabel metal5 s -8726 100906 592650 101526 6 vssa2
port 555 nsew
rlabel metal5 s -8726 64906 592650 65526 6 vssa2
port 555 nsew
rlabel metal5 s -8726 28906 592650 29526 6 vssa2
port 555 nsew
rlabel metal4 s 567834 -7654 568454 711590 6 vssa2
port 555 nsew
rlabel metal4 s 531834 -7654 532454 711590 6 vssa2
port 555 nsew
rlabel metal4 s 495834 -7654 496454 711590 6 vssa2
port 555 nsew
rlabel metal4 s 459834 -7654 460454 711590 6 vssa2
port 555 nsew
rlabel metal4 s 423834 -7654 424454 711590 6 vssa2
port 555 nsew
rlabel metal4 s 387834 -7654 388454 711590 6 vssa2
port 555 nsew
rlabel metal4 s 351834 -7654 352454 711590 6 vssa2
port 555 nsew
rlabel metal4 s 315834 -7654 316454 711590 6 vssa2
port 555 nsew
rlabel metal4 s 279834 -7654 280454 711590 6 vssa2
port 555 nsew
rlabel metal4 s 243834 -7654 244454 711590 6 vssa2
port 555 nsew
rlabel metal4 s 207834 -7654 208454 711590 6 vssa2
port 555 nsew
rlabel metal4 s 171834 -7654 172454 711590 6 vssa2
port 555 nsew
rlabel metal4 s 135834 -7654 136454 711590 6 vssa2
port 555 nsew
rlabel metal4 s 99834 -7654 100454 711590 6 vssa2
port 555 nsew
rlabel metal4 s 63834 -7654 64454 711590 6 vssa2
port 555 nsew
rlabel metal4 s 27834 -7654 28454 711590 6 vssa2
port 555 nsew
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 555 nsew
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 555 nsew
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 555 nsew
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 555 nsew
rlabel metal5 s -8726 690586 592650 691206 6 vssd1
port 556 nsew
rlabel metal5 s -8726 654586 592650 655206 6 vssd1
port 556 nsew
rlabel metal5 s -8726 618586 592650 619206 6 vssd1
port 556 nsew
rlabel metal5 s -8726 582586 592650 583206 6 vssd1
port 556 nsew
rlabel metal5 s -8726 546586 592650 547206 6 vssd1
port 556 nsew
rlabel metal5 s -8726 510586 592650 511206 6 vssd1
port 556 nsew
rlabel metal5 s -8726 474586 592650 475206 6 vssd1
port 556 nsew
rlabel metal5 s -8726 438586 592650 439206 6 vssd1
port 556 nsew
rlabel metal5 s -8726 402586 592650 403206 6 vssd1
port 556 nsew
rlabel metal5 s -8726 366586 592650 367206 6 vssd1
port 556 nsew
rlabel metal5 s -8726 330586 592650 331206 6 vssd1
port 556 nsew
rlabel metal5 s -8726 294586 592650 295206 6 vssd1
port 556 nsew
rlabel metal5 s -8726 258586 592650 259206 6 vssd1
port 556 nsew
rlabel metal5 s -8726 222586 592650 223206 6 vssd1
port 556 nsew
rlabel metal5 s -8726 186586 592650 187206 6 vssd1
port 556 nsew
rlabel metal5 s -8726 150586 592650 151206 6 vssd1
port 556 nsew
rlabel metal5 s -8726 114586 592650 115206 6 vssd1
port 556 nsew
rlabel metal5 s -8726 78586 592650 79206 6 vssd1
port 556 nsew
rlabel metal5 s -8726 42586 592650 43206 6 vssd1
port 556 nsew
rlabel metal5 s -8726 6586 592650 7206 6 vssd1
port 556 nsew
rlabel metal4 s 581514 -7654 582134 711590 6 vssd1
port 556 nsew
rlabel metal4 s 545514 -7654 546134 711590 6 vssd1
port 556 nsew
rlabel metal4 s 509514 -7654 510134 711590 6 vssd1
port 556 nsew
rlabel metal4 s 473514 -7654 474134 711590 6 vssd1
port 556 nsew
rlabel metal4 s 437514 -7654 438134 711590 6 vssd1
port 556 nsew
rlabel metal4 s 401514 -7654 402134 711590 6 vssd1
port 556 nsew
rlabel metal4 s 365514 -7654 366134 711590 6 vssd1
port 556 nsew
rlabel metal4 s 329514 -7654 330134 711590 6 vssd1
port 556 nsew
rlabel metal4 s 293514 -7654 294134 711590 6 vssd1
port 556 nsew
rlabel metal4 s 257514 -7654 258134 711590 6 vssd1
port 556 nsew
rlabel metal4 s 221514 -7654 222134 711590 6 vssd1
port 556 nsew
rlabel metal4 s 185514 -7654 186134 711590 6 vssd1
port 556 nsew
rlabel metal4 s 149514 -7654 150134 711590 6 vssd1
port 556 nsew
rlabel metal4 s 113514 -7654 114134 711590 6 vssd1
port 556 nsew
rlabel metal4 s 77514 -7654 78134 711590 6 vssd1
port 556 nsew
rlabel metal4 s 41514 -7654 42134 711590 6 vssd1
port 556 nsew
rlabel metal4 s 5514 -7654 6134 711590 6 vssd1
port 556 nsew
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 556 nsew
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 556 nsew
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 556 nsew
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 556 nsew
rlabel metal5 s -8726 698026 592650 698646 6 vssd2
port 557 nsew
rlabel metal5 s -8726 662026 592650 662646 6 vssd2
port 557 nsew
rlabel metal5 s -8726 626026 592650 626646 6 vssd2
port 557 nsew
rlabel metal5 s -8726 590026 592650 590646 6 vssd2
port 557 nsew
rlabel metal5 s -8726 554026 592650 554646 6 vssd2
port 557 nsew
rlabel metal5 s -8726 518026 592650 518646 6 vssd2
port 557 nsew
rlabel metal5 s -8726 482026 592650 482646 6 vssd2
port 557 nsew
rlabel metal5 s -8726 446026 592650 446646 6 vssd2
port 557 nsew
rlabel metal5 s -8726 410026 592650 410646 6 vssd2
port 557 nsew
rlabel metal5 s -8726 374026 592650 374646 6 vssd2
port 557 nsew
rlabel metal5 s -8726 338026 592650 338646 6 vssd2
port 557 nsew
rlabel metal5 s -8726 302026 592650 302646 6 vssd2
port 557 nsew
rlabel metal5 s -8726 266026 592650 266646 6 vssd2
port 557 nsew
rlabel metal5 s -8726 230026 592650 230646 6 vssd2
port 557 nsew
rlabel metal5 s -8726 194026 592650 194646 6 vssd2
port 557 nsew
rlabel metal5 s -8726 158026 592650 158646 6 vssd2
port 557 nsew
rlabel metal5 s -8726 122026 592650 122646 6 vssd2
port 557 nsew
rlabel metal5 s -8726 86026 592650 86646 6 vssd2
port 557 nsew
rlabel metal5 s -8726 50026 592650 50646 6 vssd2
port 557 nsew
rlabel metal5 s -8726 14026 592650 14646 6 vssd2
port 557 nsew
rlabel metal4 s 552954 -7654 553574 711590 6 vssd2
port 557 nsew
rlabel metal4 s 516954 -7654 517574 711590 6 vssd2
port 557 nsew
rlabel metal4 s 480954 -7654 481574 711590 6 vssd2
port 557 nsew
rlabel metal4 s 444954 -7654 445574 711590 6 vssd2
port 557 nsew
rlabel metal4 s 408954 -7654 409574 711590 6 vssd2
port 557 nsew
rlabel metal4 s 372954 -7654 373574 711590 6 vssd2
port 557 nsew
rlabel metal4 s 336954 -7654 337574 711590 6 vssd2
port 557 nsew
rlabel metal4 s 300954 -7654 301574 711590 6 vssd2
port 557 nsew
rlabel metal4 s 264954 -7654 265574 711590 6 vssd2
port 557 nsew
rlabel metal4 s 228954 -7654 229574 711590 6 vssd2
port 557 nsew
rlabel metal4 s 192954 -7654 193574 711590 6 vssd2
port 557 nsew
rlabel metal4 s 156954 -7654 157574 711590 6 vssd2
port 557 nsew
rlabel metal4 s 120954 -7654 121574 711590 6 vssd2
port 557 nsew
rlabel metal4 s 84954 -7654 85574 711590 6 vssd2
port 557 nsew
rlabel metal4 s 48954 -7654 49574 711590 6 vssd2
port 557 nsew
rlabel metal4 s 12954 -7654 13574 711590 6 vssd2
port 557 nsew
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 557 nsew
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 557 nsew
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 557 nsew
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 557 nsew
rlabel metal3 s 583520 258348 584960 258588 6 wb_clk_i
port 558 nsew
rlabel metal3 s -960 350828 480 351068 4 wb_rst_i
port 559 nsew
rlabel metal3 s 583520 383468 584960 383708 6 wbs_ack_o
port 560 nsew
rlabel metal2 s 199630 703520 199742 704960 6 wbs_adr_i[0]
port 561 nsew
rlabel metal2 s 54730 703520 54842 704960 6 wbs_adr_i[10]
port 562 nsew
rlabel metal3 s -960 471868 480 472108 4 wbs_adr_i[11]
port 563 nsew
rlabel metal2 s 64390 -960 64502 480 8 wbs_adr_i[12]
port 564 nsew
rlabel metal2 s 389610 -960 389722 480 8 wbs_adr_i[13]
port 565 nsew
rlabel metal3 s 583520 657508 584960 657748 6 wbs_adr_i[14]
port 566 nsew
rlabel metal3 s 583520 613308 584960 613548 6 wbs_adr_i[15]
port 567 nsew
rlabel metal2 s 443062 -960 443174 480 8 wbs_adr_i[16]
port 568 nsew
rlabel metal3 s 583520 556868 584960 557108 6 wbs_adr_i[17]
port 569 nsew
rlabel metal3 s 583520 343348 584960 343588 6 wbs_adr_i[18]
port 570 nsew
rlabel metal3 s 583520 89028 584960 89268 6 wbs_adr_i[19]
port 571 nsew
rlabel metal2 s 207358 703520 207470 704960 6 wbs_adr_i[1]
port 572 nsew
rlabel metal2 s 406354 703520 406466 704960 6 wbs_adr_i[20]
port 573 nsew
rlabel metal2 s 393474 -960 393586 480 8 wbs_adr_i[21]
port 574 nsew
rlabel metal2 s 557694 -960 557806 480 8 wbs_adr_i[22]
port 575 nsew
rlabel metal3 s 583520 278748 584960 278988 6 wbs_adr_i[23]
port 576 nsew
rlabel metal3 s -960 556188 480 556428 4 wbs_adr_i[24]
port 577 nsew
rlabel metal2 s 374154 -960 374266 480 8 wbs_adr_i[25]
port 578 nsew
rlabel metal2 s 72118 -960 72230 480 8 wbs_adr_i[26]
port 579 nsew
rlabel metal3 s -960 19668 480 19908 4 wbs_adr_i[27]
port 580 nsew
rlabel metal3 s 583520 524228 584960 524468 6 wbs_adr_i[28]
port 581 nsew
rlabel metal2 s 497802 703520 497914 704960 6 wbs_adr_i[29]
port 582 nsew
rlabel metal2 s 267250 -960 267362 480 8 wbs_adr_i[2]
port 583 nsew
rlabel metal2 s 333582 703520 333694 704960 6 wbs_adr_i[30]
port 584 nsew
rlabel metal3 s 583520 403868 584960 404108 6 wbs_adr_i[31]
port 585 nsew
rlabel metal2 s 530646 -960 530758 480 8 wbs_adr_i[3]
port 586 nsew
rlabel metal2 s 321990 703520 322102 704960 6 wbs_adr_i[4]
port 587 nsew
rlabel metal3 s -960 108748 480 108988 4 wbs_adr_i[5]
port 588 nsew
rlabel metal2 s 213798 -960 213910 480 8 wbs_adr_i[6]
port 589 nsew
rlabel metal2 s 34122 -960 34234 480 8 wbs_adr_i[7]
port 590 nsew
rlabel metal3 s 583520 97188 584960 97428 6 wbs_adr_i[8]
port 591 nsew
rlabel metal3 s 583520 290308 584960 290548 6 wbs_adr_i[9]
port 592 nsew
rlabel metal2 s 31546 703520 31658 704960 6 wbs_cyc_i
port 593 nsew
rlabel metal2 s 574438 703520 574550 704960 6 wbs_dat_i[0]
port 594 nsew
rlabel metal3 s -960 358988 480 359228 4 wbs_dat_i[10]
port 595 nsew
rlabel metal3 s -960 407268 480 407508 4 wbs_dat_i[11]
port 596 nsew
rlabel metal3 s -960 390948 480 391188 4 wbs_dat_i[12]
port 597 nsew
rlabel metal2 s 26394 -960 26506 480 8 wbs_dat_i[13]
port 598 nsew
rlabel metal2 s 144890 -960 145002 480 8 wbs_dat_i[14]
port 599 nsew
rlabel metal3 s 583520 456228 584960 456468 6 wbs_dat_i[15]
port 600 nsew
rlabel metal2 s 385746 -960 385858 480 8 wbs_dat_i[16]
port 601 nsew
rlabel metal2 s 291722 703520 291834 704960 6 wbs_dat_i[17]
port 602 nsew
rlabel metal2 s 455942 703520 456054 704960 6 wbs_dat_i[18]
port 603 nsew
rlabel metal3 s -960 576588 480 576828 4 wbs_dat_i[19]
port 604 nsew
rlabel metal2 s 103030 -960 103142 480 8 wbs_dat_i[1]
port 605 nsew
rlabel metal3 s 583520 508588 584960 508828 6 wbs_dat_i[20]
port 606 nsew
rlabel metal2 s 482346 703520 482458 704960 6 wbs_dat_i[21]
port 607 nsew
rlabel metal3 s -960 265828 480 266068 4 wbs_dat_i[22]
port 608 nsew
rlabel metal3 s 583520 629628 584960 629868 6 wbs_dat_i[23]
port 609 nsew
rlabel metal3 s 583520 310708 584960 310948 6 wbs_dat_i[24]
port 610 nsew
rlabel metal2 s 457874 -960 457986 480 8 wbs_dat_i[25]
port 611 nsew
rlabel metal2 s 410218 703520 410330 704960 6 wbs_dat_i[26]
port 612 nsew
rlabel metal2 s 19954 703520 20066 704960 6 wbs_dat_i[27]
port 613 nsew
rlabel metal2 s 206070 -960 206182 480 8 wbs_dat_i[28]
port 614 nsew
rlabel metal3 s 583520 496348 584960 496588 6 wbs_dat_i[29]
port 615 nsew
rlabel metal2 s 538374 -960 538486 480 8 wbs_dat_i[2]
port 616 nsew
rlabel metal3 s 583520 282828 584960 283068 6 wbs_dat_i[30]
port 617 nsew
rlabel metal3 s -960 249508 480 249748 4 wbs_dat_i[31]
port 618 nsew
rlabel metal3 s 583520 101268 584960 101508 6 wbs_dat_i[3]
port 619 nsew
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_i[4]
port 620 nsew
rlabel metal2 s 324566 -960 324678 480 8 wbs_dat_i[5]
port 621 nsew
rlabel metal3 s -960 3348 480 3588 4 wbs_dat_i[6]
port 622 nsew
rlabel metal2 s 398626 703520 398738 704960 6 wbs_dat_i[7]
port 623 nsew
rlabel metal3 s 583520 686068 584960 686308 6 wbs_dat_i[8]
port 624 nsew
rlabel metal3 s 583520 104668 584960 104908 6 wbs_dat_i[9]
port 625 nsew
rlabel metal2 s 53442 -960 53554 480 8 wbs_dat_o[0]
port 626 nsew
rlabel metal3 s 583520 460308 584960 460548 6 wbs_dat_o[10]
port 627 nsew
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[11]
port 628 nsew
rlabel metal3 s 583520 694228 584960 694468 6 wbs_dat_o[12]
port 629 nsew
rlabel metal2 s 383170 703520 383282 704960 6 wbs_dat_o[13]
port 630 nsew
rlabel metal3 s 583520 145468 584960 145708 6 wbs_dat_o[14]
port 631 nsew
rlabel metal2 s 363850 703520 363962 704960 6 wbs_dat_o[15]
port 632 nsew
rlabel metal3 s -960 116908 480 117148 4 wbs_dat_o[16]
port 633 nsew
rlabel metal3 s -960 136628 480 136868 4 wbs_dat_o[17]
port 634 nsew
rlabel metal2 s 435334 -960 435446 480 8 wbs_dat_o[18]
port 635 nsew
rlabel metal2 s -10 -960 102 480 8 wbs_dat_o[19]
port 636 nsew
rlabel metal2 s 508106 -960 508218 480 8 wbs_dat_o[1]
port 637 nsew
rlabel metal3 s -960 257668 480 257908 4 wbs_dat_o[20]
port 638 nsew
rlabel metal3 s -960 524228 480 524468 4 wbs_dat_o[21]
port 639 nsew
rlabel metal2 s 92726 703520 92838 704960 6 wbs_dat_o[22]
port 640 nsew
rlabel metal3 s -960 169268 480 169508 4 wbs_dat_o[23]
port 641 nsew
rlabel metal2 s 133298 -960 133410 480 8 wbs_dat_o[24]
port 642 nsew
rlabel metal2 s 49578 -960 49690 480 8 wbs_dat_o[25]
port 643 nsew
rlabel metal2 s 256946 703520 257058 704960 6 wbs_dat_o[26]
port 644 nsew
rlabel metal2 s 112046 703520 112158 704960 6 wbs_dat_o[27]
port 645 nsew
rlabel metal2 s 347106 -960 347218 480 8 wbs_dat_o[28]
port 646 nsew
rlabel metal2 s 367714 703520 367826 704960 6 wbs_dat_o[29]
port 647 nsew
rlabel metal3 s 583520 242028 584960 242268 6 wbs_dat_o[2]
port 648 nsew
rlabel metal3 s -960 403188 480 403428 4 wbs_dat_o[30]
port 649 nsew
rlabel metal3 s 583520 569108 584960 569348 6 wbs_dat_o[31]
port 650 nsew
rlabel metal2 s 141026 -960 141138 480 8 wbs_dat_o[3]
port 651 nsew
rlabel metal2 s 244066 -960 244178 480 8 wbs_dat_o[4]
port 652 nsew
rlabel metal3 s -960 35988 480 36228 4 wbs_dat_o[5]
port 653 nsew
rlabel metal3 s 583520 544628 584960 544868 6 wbs_dat_o[6]
port 654 nsew
rlabel metal2 s 381882 -960 381994 480 8 wbs_dat_o[7]
port 655 nsew
rlabel metal2 s 359986 703520 360098 704960 6 wbs_dat_o[8]
port 656 nsew
rlabel metal2 s 352902 703520 353014 704960 6 wbs_dat_o[9]
port 657 nsew
rlabel metal3 s -960 600388 480 600628 4 wbs_sel_i[0]
port 658 nsew
rlabel metal2 s 16090 703520 16202 704960 6 wbs_sel_i[1]
port 659 nsew
rlabel metal2 s 454654 -960 454766 480 8 wbs_sel_i[2]
port 660 nsew
rlabel metal3 s -960 140708 480 140948 4 wbs_sel_i[3]
port 661 nsew
rlabel metal3 s -960 543948 480 544188 4 wbs_stb_i
port 662 nsew
rlabel metal3 s 583520 371228 584960 371468 6 wbs_we_i
port 663 nsew
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 139800590
string GDS_FILE /home/passant/caravel_user_project_analog/openlane/user_analog_project_wrapper/runs/23_05_22_01_01/results/signoff/user_analog_project_wrapper.magic.gds
string GDS_START 135332
<< end >>

