VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_analog_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_analog_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN gpio_analog[0]
    PORT
      LAYER met2 ;
        RECT 437.870 -4.800 438.430 2.400 ;
    END
  END gpio_analog[0]
  PIN gpio_analog[10]
    PORT
      LAYER met2 ;
        RECT 782.410 -4.800 782.970 2.400 ;
    END
  END gpio_analog[10]
  PIN gpio_analog[11]
    PORT
      LAYER met3 ;
        RECT 2917.600 281.940 2924.800 283.140 ;
    END
  END gpio_analog[11]
  PIN gpio_analog[12]
    PORT
      LAYER met2 ;
        RECT 502.270 3517.600 502.830 3524.800 ;
    END
  END gpio_analog[12]
  PIN gpio_analog[13]
    PORT
      LAYER met3 ;
        RECT -4.800 1631.740 2.400 1632.940 ;
    END
  END gpio_analog[13]
  PIN gpio_analog[14]
    PORT
      LAYER met2 ;
        RECT 1725.870 3517.600 1726.430 3524.800 ;
    END
  END gpio_analog[14]
  PIN gpio_analog[15]
    PORT
      LAYER met3 ;
        RECT 2917.600 1111.540 2924.800 1112.740 ;
    END
  END gpio_analog[15]
  PIN gpio_analog[16]
    PORT
      LAYER met3 ;
        RECT -4.800 3185.540 2.400 3186.740 ;
    END
  END gpio_analog[16]
  PIN gpio_analog[17]
    PORT
      LAYER met3 ;
        RECT -4.800 642.340 2.400 643.540 ;
    END
  END gpio_analog[17]
  PIN gpio_analog[1]
    PORT
      LAYER met3 ;
        RECT 2917.600 404.340 2924.800 405.540 ;
    END
  END gpio_analog[1]
  PIN gpio_analog[2]
    PORT
      LAYER met2 ;
        RECT 1297.610 -4.800 1298.170 2.400 ;
    END
  END gpio_analog[2]
  PIN gpio_analog[3]
    PORT
      LAYER met3 ;
        RECT -4.800 2175.740 2.400 2176.940 ;
    END
  END gpio_analog[3]
  PIN gpio_analog[4]
    PORT
      LAYER met3 ;
        RECT 2917.600 3369.140 2924.800 3370.340 ;
    END
  END gpio_analog[4]
  PIN gpio_analog[5]
    PORT
      LAYER met3 ;
        RECT -4.800 1026.540 2.400 1027.740 ;
    END
  END gpio_analog[5]
  PIN gpio_analog[6]
    PORT
      LAYER met3 ;
        RECT -4.800 1995.540 2.400 1996.740 ;
    END
  END gpio_analog[6]
  PIN gpio_analog[7]
    PORT
      LAYER met2 ;
        RECT 379.910 -4.800 380.470 2.400 ;
    END
  END gpio_analog[7]
  PIN gpio_analog[8]
    PORT
      LAYER met2 ;
        RECT 2730.510 -4.800 2731.070 2.400 ;
    END
  END gpio_analog[8]
  PIN gpio_analog[9]
    PORT
      LAYER met2 ;
        RECT 2060.750 -4.800 2061.310 2.400 ;
    END
  END gpio_analog[9]
  PIN gpio_noesd[0]
    PORT
      LAYER met2 ;
        RECT 1201.010 -4.800 1201.570 2.400 ;
    END
  END gpio_noesd[0]
  PIN gpio_noesd[10]
    PORT
      LAYER met3 ;
        RECT -4.800 2682.340 2.400 2683.540 ;
    END
  END gpio_noesd[10]
  PIN gpio_noesd[11]
    PORT
      LAYER met3 ;
        RECT -4.800 2236.940 2.400 2238.140 ;
    END
  END gpio_noesd[11]
  PIN gpio_noesd[12]
    PORT
      LAYER met2 ;
        RECT 866.130 3517.600 866.690 3524.800 ;
    END
  END gpio_noesd[12]
  PIN gpio_noesd[13]
    PORT
      LAYER met2 ;
        RECT 1954.490 3517.600 1955.050 3524.800 ;
    END
  END gpio_noesd[13]
  PIN gpio_noesd[14]
    PORT
      LAYER met3 ;
        RECT -4.800 1913.940 2.400 1915.140 ;
    END
  END gpio_noesd[14]
  PIN gpio_noesd[15]
    PORT
      LAYER met3 ;
        RECT -4.800 298.940 2.400 300.140 ;
    END
  END gpio_noesd[15]
  PIN gpio_noesd[16]
    PORT
      LAYER met3 ;
        RECT 2917.600 142.540 2924.800 143.740 ;
    END
  END gpio_noesd[16]
  PIN gpio_noesd[17]
    PORT
      LAYER met2 ;
        RECT 1056.110 3517.600 1056.670 3524.800 ;
    END
  END gpio_noesd[17]
  PIN gpio_noesd[1]
    PORT
      LAYER met2 ;
        RECT 608.530 -4.800 609.090 2.400 ;
    END
  END gpio_noesd[1]
  PIN gpio_noesd[2]
    PORT
      LAYER met2 ;
        RECT 1642.150 -4.800 1642.710 2.400 ;
    END
  END gpio_noesd[2]
  PIN gpio_noesd[3]
    PORT
      LAYER met3 ;
        RECT 2917.600 3209.340 2924.800 3210.540 ;
    END
  END gpio_noesd[3]
  PIN gpio_noesd[4]
    PORT
      LAYER met2 ;
        RECT 959.510 3517.600 960.070 3524.800 ;
    END
  END gpio_noesd[4]
  PIN gpio_noesd[5]
    PORT
      LAYER met3 ;
        RECT 2917.600 322.740 2924.800 323.940 ;
    END
  END gpio_noesd[5]
  PIN gpio_noesd[6]
    PORT
      LAYER met3 ;
        RECT 2917.600 3005.340 2924.800 3006.540 ;
    END
  END gpio_noesd[6]
  PIN gpio_noesd[7]
    PORT
      LAYER met3 ;
        RECT 2917.600 2461.340 2924.800 2462.540 ;
    END
  END gpio_noesd[7]
  PIN gpio_noesd[8]
    PORT
      LAYER met3 ;
        RECT -4.800 441.740 2.400 442.940 ;
    END
  END gpio_noesd[8]
  PIN gpio_noesd[9]
    PORT
      LAYER met3 ;
        RECT -4.800 662.740 2.400 663.940 ;
    END
  END gpio_noesd[9]
  PIN io_analog[0]
    PORT
      LAYER met3 ;
        RECT -4.800 1227.140 2.400 1228.340 ;
    END
  END io_analog[0]
  PIN io_analog[10]
    PORT
      LAYER met2 ;
        RECT 283.310 -4.800 283.870 2.400 ;
    END
  END io_analog[10]
  PIN io_analog[1]
    PORT
      LAYER met3 ;
        RECT 2917.600 302.340 2924.800 303.540 ;
    END
  END io_analog[1]
  PIN io_analog[2]
    PORT
      LAYER met3 ;
        RECT 2917.600 2763.940 2924.800 2765.140 ;
    END
  END io_analog[2]
  PIN io_analog[3]
    PORT
      LAYER met2 ;
        RECT 1143.050 -4.800 1143.610 2.400 ;
    END
  END io_analog[3]
  PIN io_analog[4]
    PORT
      LAYER met2 ;
        RECT 569.890 -4.800 570.450 2.400 ;
    END
  END io_analog[4]
  PIN io_analog[5]
    PORT
      LAYER met2 ;
        RECT 444.310 3517.600 444.870 3524.800 ;
    END
  END io_analog[5]
  PIN io_analog[6]
    PORT
      LAYER met2 ;
        RECT 2253.950 -4.800 2254.510 2.400 ;
    END
  END io_analog[6]
  PIN io_analog[7]
    PORT
      LAYER met3 ;
        RECT -4.800 1169.340 2.400 1170.540 ;
    END
  END io_analog[7]
  PIN io_analog[8]
    PORT
      LAYER met2 ;
        RECT 1049.670 -4.800 1050.230 2.400 ;
    END
  END io_analog[8]
  PIN io_analog[9]
    PORT
      LAYER met3 ;
        RECT -4.800 1672.540 2.400 1673.740 ;
    END
  END io_analog[9]
  PIN io_clamp_high[0]
    PORT
      LAYER met2 ;
        RECT 112.650 -4.800 113.210 2.400 ;
    END
  END io_clamp_high[0]
  PIN io_clamp_high[1]
    PORT
      LAYER met3 ;
        RECT 2917.600 2906.740 2924.800 2907.940 ;
    END
  END io_clamp_high[1]
  PIN io_clamp_high[2]
    PORT
      LAYER met3 ;
        RECT 2917.600 1815.340 2924.800 1816.540 ;
    END
  END io_clamp_high[2]
  PIN io_clamp_low[0]
    PORT
      LAYER met3 ;
        RECT -4.800 621.940 2.400 623.140 ;
    END
  END io_clamp_low[0]
  PIN io_clamp_low[1]
    PORT
      LAYER met2 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END io_clamp_low[1]
  PIN io_clamp_low[2]
    PORT
      LAYER met3 ;
        RECT -4.800 3246.740 2.400 3247.940 ;
    END
  END io_clamp_low[2]
  PIN io_in[0]
    PORT
      LAYER met2 ;
        RECT 189.930 -4.800 190.490 2.400 ;
    END
  END io_in[0]
  PIN io_in[10]
    PORT
      LAYER met3 ;
        RECT 2917.600 2522.540 2924.800 2523.740 ;
    END
  END io_in[10]
  PIN io_in[11]
    PORT
      LAYER met2 ;
        RECT 2469.690 3517.600 2470.250 3524.800 ;
    END
  END io_in[11]
  PIN io_in[12]
    PORT
      LAYER met2 ;
        RECT 2012.450 3517.600 2013.010 3524.800 ;
    END
  END io_in[12]
  PIN io_in[13]
    PORT
      LAYER met2 ;
        RECT 495.830 -4.800 496.390 2.400 ;
    END
  END io_in[13]
  PIN io_in[14]
    PORT
      LAYER met2 ;
        RECT 2080.070 -4.800 2080.630 2.400 ;
    END
  END io_in[14]
  PIN io_in[15]
    PORT
      LAYER met3 ;
        RECT -4.800 380.540 2.400 381.740 ;
    END
  END io_in[15]
  PIN io_in[16]
    PORT
      LAYER met2 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END io_in[16]
  PIN io_in[17]
    PORT
      LAYER met3 ;
        RECT 2917.600 1189.740 2924.800 1190.940 ;
    END
  END io_in[17]
  PIN io_in[18]
    PORT
      LAYER met3 ;
        RECT 2917.600 363.540 2924.800 364.740 ;
    END
  END io_in[18]
  PIN io_in[19]
    PORT
      LAYER met3 ;
        RECT -4.800 2821.740 2.400 2822.940 ;
    END
  END io_in[19]
  PIN io_in[1]
    PORT
      LAYER met2 ;
        RECT 2463.250 -4.800 2463.810 2.400 ;
    END
  END io_in[1]
  PIN io_in[20]
    PORT
      LAYER met2 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END io_in[20]
  PIN io_in[21]
    PORT
      LAYER met2 ;
        RECT 1680.790 -4.800 1681.350 2.400 ;
    END
  END io_in[21]
  PIN io_in[22]
    PORT
      LAYER met3 ;
        RECT 2917.600 666.140 2924.800 667.340 ;
    END
  END io_in[22]
  PIN io_in[23]
    PORT
      LAYER met2 ;
        RECT 1323.370 3517.600 1323.930 3524.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    PORT
      LAYER met3 ;
        RECT 2917.600 1998.940 2924.800 2000.140 ;
    END
  END io_in[24]
  PIN io_in[25]
    PORT
      LAYER met2 ;
        RECT 2901.170 -4.800 2901.730 2.400 ;
    END
  END io_in[25]
  PIN io_in[26]
    PORT
      LAYER met2 ;
        RECT 2678.990 3517.600 2679.550 3524.800 ;
    END
  END io_in[26]
  PIN io_in[2]
    PORT
      LAYER met3 ;
        RECT 2917.600 2260.740 2924.800 2261.940 ;
    END
  END io_in[2]
  PIN io_in[3]
    PORT
      LAYER met3 ;
        RECT -4.800 1570.540 2.400 1571.740 ;
    END
  END io_in[3]
  PIN io_in[4]
    PORT
      LAYER met2 ;
        RECT 2138.030 -4.800 2138.590 2.400 ;
    END
  END io_in[4]
  PIN io_in[5]
    PORT
      LAYER met2 ;
        RECT 653.610 3517.600 654.170 3524.800 ;
    END
  END io_in[5]
  PIN io_in[6]
    PORT
      LAYER met3 ;
        RECT 2917.600 2743.540 2924.800 2744.740 ;
    END
  END io_in[6]
  PIN io_in[7]
    PORT
      LAYER met3 ;
        RECT -4.800 281.940 2.400 283.140 ;
    END
  END io_in[7]
  PIN io_in[8]
    PORT
      LAYER met2 ;
        RECT 418.550 -4.800 419.110 2.400 ;
    END
  END io_in[8]
  PIN io_in[9]
    PORT
      LAYER met2 ;
        RECT 1152.710 3517.600 1153.270 3524.800 ;
    END
  END io_in[9]
  PIN io_in_3v3[0]
    PORT
      LAYER met2 ;
        RECT 821.050 -4.800 821.610 2.400 ;
    END
  END io_in_3v3[0]
  PIN io_in_3v3[10]
    PORT
      LAYER met2 ;
        RECT 228.570 -4.800 229.130 2.400 ;
    END
  END io_in_3v3[10]
  PIN io_in_3v3[11]
    PORT
      LAYER met2 ;
        RECT 1687.230 3517.600 1687.790 3524.800 ;
    END
  END io_in_3v3[11]
  PIN io_in_3v3[12]
    PORT
      LAYER met2 ;
        RECT 2659.670 3517.600 2660.230 3524.800 ;
    END
  END io_in_3v3[12]
  PIN io_in_3v3[13]
    PORT
      LAYER met2 ;
        RECT 54.690 -4.800 55.250 2.400 ;
    END
  END io_in_3v3[13]
  PIN io_in_3v3[14]
    PORT
      LAYER met3 ;
        RECT -4.800 3205.940 2.400 3207.140 ;
    END
  END io_in_3v3[14]
  PIN io_in_3v3[15]
    PORT
      LAYER met3 ;
        RECT 2917.600 1029.940 2924.800 1031.140 ;
    END
  END io_in_3v3[15]
  PIN io_in_3v3[16]
    PORT
      LAYER met3 ;
        RECT 2917.600 788.540 2924.800 789.740 ;
    END
  END io_in_3v3[16]
  PIN io_in_3v3[17]
    PORT
      LAYER met3 ;
        RECT -4.800 3287.540 2.400 3288.740 ;
    END
  END io_in_3v3[17]
  PIN io_in_3v3[18]
    PORT
      LAYER met3 ;
        RECT -4.800 1832.340 2.400 1833.540 ;
    END
  END io_in_3v3[18]
  PIN io_in_3v3[19]
    PORT
      LAYER met3 ;
        RECT -4.800 3165.140 2.400 3166.340 ;
    END
  END io_in_3v3[19]
  PIN io_in_3v3[1]
    PORT
      LAYER met3 ;
        RECT 2917.600 261.540 2924.800 262.740 ;
    END
  END io_in_3v3[1]
  PIN io_in_3v3[20]
    PORT
      LAYER met2 ;
        RECT 367.030 3517.600 367.590 3524.800 ;
    END
  END io_in_3v3[20]
  PIN io_in_3v3[21]
    PORT
      LAYER met3 ;
        RECT -4.800 2964.540 2.400 2965.740 ;
    END
  END io_in_3v3[21]
  PIN io_in_3v3[22]
    PORT
      LAYER met3 ;
        RECT -4.800 3488.140 2.400 3489.340 ;
    END
  END io_in_3v3[22]
  PIN io_in_3v3[23]
    PORT
      LAYER met3 ;
        RECT -4.800 3386.140 2.400 3387.340 ;
    END
  END io_in_3v3[23]
  PIN io_in_3v3[24]
    PORT
      LAYER met2 ;
        RECT 1468.270 -4.800 1468.830 2.400 ;
    END
  END io_in_3v3[24]
  PIN io_in_3v3[25]
    PORT
      LAYER met3 ;
        RECT 2917.600 1675.940 2924.800 1677.140 ;
    END
  END io_in_3v3[25]
  PIN io_in_3v3[26]
    PORT
      LAYER met3 ;
        RECT -4.800 1975.140 2.400 1976.340 ;
    END
  END io_in_3v3[26]
  PIN io_in_3v3[2]
    PORT
      LAYER met2 ;
        RECT 6.390 3517.600 6.950 3524.800 ;
    END
  END io_in_3v3[2]
  PIN io_in_3v3[3]
    PORT
      LAYER met3 ;
        RECT 2917.600 3267.140 2924.800 3268.340 ;
    END
  END io_in_3v3[3]
  PIN io_in_3v3[4]
    PORT
      LAYER met2 ;
        RECT 2833.550 3517.600 2834.110 3524.800 ;
    END
  END io_in_3v3[4]
  PIN io_in_3v3[5]
    PORT
      LAYER met2 ;
        RECT 1564.870 -4.800 1565.430 2.400 ;
    END
  END io_in_3v3[5]
  PIN io_in_3v3[6]
    PORT
      LAYER met2 ;
        RECT 2234.630 -4.800 2235.190 2.400 ;
    END
  END io_in_3v3[6]
  PIN io_in_3v3[7]
    PORT
      LAYER met2 ;
        RECT 991.710 -4.800 992.270 2.400 ;
    END
  END io_in_3v3[7]
  PIN io_in_3v3[8]
    PORT
      LAYER met2 ;
        RECT 1477.930 3517.600 1478.490 3524.800 ;
    END
  END io_in_3v3[8]
  PIN io_in_3v3[9]
    PORT
      LAYER met2 ;
        RECT 2769.150 -4.800 2769.710 2.400 ;
    END
  END io_in_3v3[9]
  PIN io_oeb[0]
    PORT
      LAYER met3 ;
        RECT -4.800 2379.740 2.400 2380.940 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    PORT
      LAYER met2 ;
        RECT 2373.090 3517.600 2373.650 3524.800 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    PORT
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    PORT
      LAYER met2 ;
        RECT 1832.130 -4.800 1832.690 2.400 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    PORT
      LAYER met2 ;
        RECT 2575.950 -4.800 2576.510 2.400 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    PORT
      LAYER met3 ;
        RECT 2917.600 1754.140 2924.800 1755.340 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    PORT
      LAYER met3 ;
        RECT -4.800 2437.540 2.400 2438.740 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    PORT
      LAYER met3 ;
        RECT -4.800 2641.540 2.400 2642.740 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    PORT
      LAYER met3 ;
        RECT 2917.600 2964.540 2924.800 2965.740 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    PORT
      LAYER met2 ;
        RECT 647.170 -4.800 647.730 2.400 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    PORT
      LAYER met3 ;
        RECT 2917.600 3246.740 2924.800 3247.940 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    PORT
      LAYER met2 ;
        RECT 2508.330 3517.600 2508.890 3524.800 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    PORT
      LAYER met2 ;
        RECT 2624.250 3517.600 2624.810 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    PORT
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    PORT
      LAYER met2 ;
        RECT 302.630 -4.800 303.190 2.400 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    PORT
      LAYER met3 ;
        RECT 2917.600 846.340 2924.800 847.540 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    PORT
      LAYER met2 ;
        RECT 1745.190 3517.600 1745.750 3524.800 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    PORT
      LAYER met3 ;
        RECT 2917.600 2420.540 2924.800 2421.740 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    PORT
      LAYER met3 ;
        RECT 2917.600 1876.540 2924.800 1877.740 ;
    END
  END io_oeb[26]
  PIN io_oeb[2]
    PORT
      LAYER met3 ;
        RECT -4.800 3042.740 2.400 3043.940 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    PORT
      LAYER met3 ;
        RECT -4.800 3124.340 2.400 3125.540 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    PORT
      LAYER met3 ;
        RECT -4.800 2338.940 2.400 2340.140 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    PORT
      LAYER met3 ;
        RECT 2917.600 2804.740 2924.800 2805.940 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    PORT
      LAYER met2 ;
        RECT 196.370 3517.600 196.930 3524.800 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    PORT
      LAYER met3 ;
        RECT -4.800 2600.740 2.400 2601.940 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    PORT
      LAYER met2 ;
        RECT 1497.250 3517.600 1497.810 3524.800 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    PORT
      LAYER met3 ;
        RECT 2917.600 1471.940 2924.800 1473.140 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    PORT
      LAYER met2 ;
        RECT 2604.930 3517.600 2605.490 3524.800 ;
    END
  END io_out[0]
  PIN io_out[10]
    PORT
      LAYER met3 ;
        RECT -4.800 887.140 2.400 888.340 ;
    END
  END io_out[10]
  PIN io_out[11]
    PORT
      LAYER met3 ;
        RECT 2917.600 3328.340 2924.800 3329.540 ;
    END
  END io_out[11]
  PIN io_out[12]
    PORT
      LAYER met3 ;
        RECT -4.800 1492.340 2.400 1493.540 ;
    END
  END io_out[12]
  PIN io_out[13]
    PORT
      LAYER met3 ;
        RECT 2917.600 2077.140 2924.800 2078.340 ;
    END
  END io_out[13]
  PIN io_out[14]
    PORT
      LAYER met2 ;
        RECT 1342.690 3517.600 1343.250 3524.800 ;
    END
  END io_out[14]
  PIN io_out[15]
    PORT
      LAYER met3 ;
        RECT -4.800 1733.740 2.400 1734.940 ;
    END
  END io_out[15]
  PIN io_out[16]
    PORT
      LAYER met2 ;
        RECT 292.970 3517.600 293.530 3524.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    PORT
      LAYER met2 ;
        RECT 978.830 3517.600 979.390 3524.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    PORT
      LAYER met2 ;
        RECT 119.090 3517.600 119.650 3524.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    PORT
      LAYER met3 ;
        RECT 2917.600 1332.540 2924.800 1333.740 ;
    END
  END io_out[19]
  PIN io_out[1]
    PORT
      LAYER met3 ;
        RECT 2917.600 2036.340 2924.800 2037.540 ;
    END
  END io_out[1]
  PIN io_out[20]
    PORT
      LAYER met2 ;
        RECT 350.930 3517.600 351.490 3524.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    PORT
      LAYER met2 ;
        RECT 1355.570 -4.800 1356.130 2.400 ;
    END
  END io_out[21]
  PIN io_out[22]
    PORT
      LAYER met3 ;
        RECT -4.800 924.540 2.400 925.740 ;
    END
  END io_out[22]
  PIN io_out[23]
    PORT
      LAYER met3 ;
        RECT 2917.600 1774.540 2924.800 1775.740 ;
    END
  END io_out[23]
  PIN io_out[24]
    PORT
      LAYER met3 ;
        RECT -4.800 3426.940 2.400 3428.140 ;
    END
  END io_out[24]
  PIN io_out[25]
    PORT
      LAYER met3 ;
        RECT -4.800 1349.540 2.400 1350.740 ;
    END
  END io_out[25]
  PIN io_out[26]
    PORT
      LAYER met2 ;
        RECT 1107.630 -4.800 1108.190 2.400 ;
    END
  END io_out[26]
  PIN io_out[2]
    PORT
      LAYER met2 ;
        RECT 895.110 -4.800 895.670 2.400 ;
    END
  END io_out[2]
  PIN io_out[3]
    PORT
      LAYER met2 ;
        RECT 1381.330 3517.600 1381.890 3524.800 ;
    END
  END io_out[3]
  PIN io_out[4]
    PORT
      LAYER met2 ;
        RECT 2353.770 3517.600 2354.330 3524.800 ;
    END
  END io_out[4]
  PIN io_out[5]
    PORT
      LAYER met3 ;
        RECT -4.800 2417.140 2.400 2418.340 ;
    END
  END io_out[5]
  PIN io_out[6]
    PORT
      LAYER met3 ;
        RECT 2917.600 825.940 2924.800 827.140 ;
    END
  END io_out[6]
  PIN io_out[7]
    PORT
      LAYER met3 ;
        RECT -4.800 3267.140 2.400 3268.340 ;
    END
  END io_out[7]
  PIN io_out[8]
    PORT
      LAYER met3 ;
        RECT 2917.600 604.940 2924.800 606.140 ;
    END
  END io_out[8]
  PIN io_out[9]
    PORT
      LAYER met3 ;
        RECT 2917.600 1250.940 2924.800 1252.140 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    PORT
      LAYER met2 ;
        RECT 788.850 3517.600 789.410 3524.800 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    PORT
      LAYER met3 ;
        RECT 2917.600 3127.740 2924.800 3128.940 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    PORT
      LAYER met3 ;
        RECT 2917.600 1070.740 2924.800 1071.940 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    PORT
      LAYER met2 ;
        RECT 1935.170 3517.600 1935.730 3524.800 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    PORT
      LAYER met3 ;
        RECT 2917.600 101.740 2924.800 102.940 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    PORT
      LAYER met3 ;
        RECT -4.800 1852.740 2.400 1853.940 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    PORT
      LAYER met2 ;
        RECT 1114.070 3517.600 1114.630 3524.800 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    PORT
      LAYER met2 ;
        RECT 672.930 3517.600 673.490 3524.800 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    PORT
      LAYER met3 ;
        RECT -4.800 2077.140 2.400 2078.340 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    PORT
      LAYER met3 ;
        RECT 2917.600 2923.740 2924.800 2924.940 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    PORT
      LAYER met3 ;
        RECT -4.800 805.540 2.400 806.740 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    PORT
      LAYER met3 ;
        RECT 2917.600 1896.940 2924.800 1898.140 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    PORT
      LAYER met3 ;
        RECT -4.800 1431.140 2.400 1432.340 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    PORT
      LAYER met3 ;
        RECT 2917.600 1352.940 2924.800 1354.140 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    PORT
      LAYER met3 ;
        RECT -4.800 1873.140 2.400 1874.340 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    PORT
      LAYER met3 ;
        RECT -4.800 3365.740 2.400 3366.940 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    PORT
      LAYER met3 ;
        RECT -4.800 2580.340 2.400 2581.540 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    PORT
      LAYER met2 ;
        RECT 1629.270 3517.600 1629.830 3524.800 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    PORT
      LAYER met2 ;
        RECT 2633.910 -4.800 2634.470 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    PORT
      LAYER met3 ;
        RECT -4.800 1692.940 2.400 1694.140 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    PORT
      LAYER met3 ;
        RECT 2917.600 2604.140 2924.800 2605.340 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    PORT
      LAYER met3 ;
        RECT 2917.600 1050.340 2924.800 1051.540 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    PORT
      LAYER met2 ;
        RECT 482.950 3517.600 483.510 3524.800 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    PORT
      LAYER met3 ;
        RECT -4.800 1529.740 2.400 1530.940 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    PORT
      LAYER met2 ;
        RECT 801.730 -4.800 802.290 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    PORT
      LAYER met2 ;
        RECT 685.810 -4.800 686.370 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    PORT
      LAYER met3 ;
        RECT -4.800 2134.940 2.400 2136.140 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    PORT
      LAYER met2 ;
        RECT 2067.190 3517.600 2067.750 3524.800 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    PORT
      LAYER met2 ;
        RECT 2424.610 -4.800 2425.170 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    PORT
      LAYER met3 ;
        RECT -4.800 2097.540 2.400 2098.740 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    PORT
      LAYER met2 ;
        RECT 2794.910 3517.600 2795.470 3524.800 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    PORT
      LAYER met3 ;
        RECT 2917.600 927.940 2924.800 929.140 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    PORT
      LAYER met3 ;
        RECT 2917.600 1696.340 2924.800 1697.540 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    PORT
      LAYER met3 ;
        RECT -4.800 2699.340 2.400 2700.540 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    PORT
      LAYER met3 ;
        RECT -4.800 2740.140 2.400 2741.340 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    PORT
      LAYER met3 ;
        RECT -4.800 339.740 2.400 340.940 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    PORT
      LAYER met3 ;
        RECT -4.800 785.140 2.400 786.340 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    PORT
      LAYER met3 ;
        RECT -4.800 2257.340 2.400 2258.540 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    PORT
      LAYER met2 ;
        RECT 2241.070 3517.600 2241.630 3524.800 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    PORT
      LAYER met2 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    PORT
      LAYER met3 ;
        RECT -4.800 1550.140 2.400 1551.340 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    PORT
      LAYER met2 ;
        RECT 138.410 3517.600 138.970 3524.800 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    PORT
      LAYER met2 ;
        RECT 904.770 3517.600 905.330 3524.800 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    PORT
      LAYER met3 ;
        RECT -4.800 2196.140 2.400 2197.340 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    PORT
      LAYER met3 ;
        RECT 2917.600 2117.940 2924.800 2119.140 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    PORT
      LAYER met2 ;
        RECT 2163.790 3517.600 2164.350 3524.800 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    PORT
      LAYER met2 ;
        RECT 2521.210 -4.800 2521.770 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    PORT
      LAYER met2 ;
        RECT 1448.950 -4.800 1449.510 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    PORT
      LAYER met3 ;
        RECT -4.800 2318.540 2.400 2319.740 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    PORT
      LAYER met3 ;
        RECT -4.800 1713.340 2.400 1714.540 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    PORT
      LAYER met2 ;
        RECT 2195.990 -4.800 2196.550 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    PORT
      LAYER met3 ;
        RECT -4.800 2457.940 2.400 2459.140 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    PORT
      LAYER met3 ;
        RECT 2917.600 3025.740 2924.800 3026.940 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    PORT
      LAYER met2 ;
        RECT 1513.350 3517.600 1513.910 3524.800 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    PORT
      LAYER met3 ;
        RECT 2917.600 2944.140 2924.800 2945.340 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    PORT
      LAYER met3 ;
        RECT -4.800 37.140 2.400 38.340 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    PORT
      LAYER met3 ;
        RECT -4.800 3324.940 2.400 3326.140 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    PORT
      LAYER met2 ;
        RECT 2756.270 3517.600 2756.830 3524.800 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    PORT
      LAYER met2 ;
        RECT 2717.630 3517.600 2718.190 3524.800 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    PORT
      LAYER met2 ;
        RECT 1648.590 3517.600 1649.150 3524.800 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    PORT
      LAYER met2 ;
        RECT 743.770 -4.800 744.330 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    PORT
      LAYER met3 ;
        RECT 2917.600 1978.540 2924.800 1979.740 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    PORT
      LAYER met2 ;
        RECT 692.250 3517.600 692.810 3524.800 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    PORT
      LAYER met3 ;
        RECT -4.800 3103.940 2.400 3105.140 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    PORT
      LAYER met3 ;
        RECT -4.800 723.940 2.400 725.140 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    PORT
      LAYER met3 ;
        RECT 2917.600 1594.340 2924.800 1595.540 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    PORT
      LAYER met3 ;
        RECT -4.800 2298.140 2.400 2299.340 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    PORT
      LAYER met2 ;
        RECT 405.670 3517.600 406.230 3524.800 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    PORT
      LAYER met2 ;
        RECT 618.190 3517.600 618.750 3524.800 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    PORT
      LAYER met3 ;
        RECT -4.800 2903.340 2.400 2904.540 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    PORT
      LAYER met3 ;
        RECT 2917.600 2097.540 2924.800 2098.740 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    PORT
      LAYER met3 ;
        RECT 2917.600 162.940 2924.800 164.140 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    PORT
      LAYER met2 ;
        RECT 2157.350 -4.800 2157.910 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    PORT
      LAYER met2 ;
        RECT 2443.930 -4.800 2444.490 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    PORT
      LAYER met3 ;
        RECT 2917.600 2502.140 2924.800 2503.340 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    PORT
      LAYER met3 ;
        RECT -4.800 2760.540 2.400 2761.740 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    PORT
      LAYER met2 ;
        RECT 1278.290 -4.800 1278.850 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    PORT
      LAYER met2 ;
        RECT 16.050 -4.800 16.610 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    PORT
      LAYER met3 ;
        RECT 2917.600 1614.740 2924.800 1615.940 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    PORT
      LAYER met3 ;
        RECT -4.800 2539.540 2.400 2540.740 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    PORT
      LAYER met3 ;
        RECT 2917.600 2056.740 2924.800 2057.940 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    PORT
      LAYER met2 ;
        RECT 1973.810 3517.600 1974.370 3524.800 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    PORT
      LAYER met3 ;
        RECT -4.800 523.340 2.400 524.540 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    PORT
      LAYER met3 ;
        RECT -4.800 3063.140 2.400 3064.340 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    PORT
      LAYER met2 ;
        RECT 2711.190 -4.800 2711.750 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    PORT
      LAYER met2 ;
        RECT 2843.210 -4.800 2843.770 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    PORT
      LAYER met3 ;
        RECT 2917.600 241.140 2924.800 242.340 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    PORT
      LAYER met3 ;
        RECT -4.800 944.940 2.400 946.140 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    PORT
      LAYER met3 ;
        RECT 2917.600 866.740 2924.800 867.940 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    PORT
      LAYER met3 ;
        RECT 2917.600 2886.340 2924.800 2887.540 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    PORT
      LAYER met3 ;
        RECT 2917.600 1655.540 2924.800 1656.740 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    PORT
      LAYER met2 ;
        RECT 399.230 -4.800 399.790 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    PORT
      LAYER met3 ;
        RECT 2917.600 2825.140 2924.800 2826.340 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    PORT
      LAYER met3 ;
        RECT 2917.600 3389.540 2924.800 3390.740 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    PORT
      LAYER met3 ;
        RECT 2917.600 1492.340 2924.800 1493.540 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    PORT
      LAYER met3 ;
        RECT -4.800 2498.740 2.400 2499.940 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    PORT
      LAYER met3 ;
        RECT -4.800 825.940 2.400 827.140 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    PORT
      LAYER met2 ;
        RECT 312.290 3517.600 312.850 3524.800 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    PORT
      LAYER met3 ;
        RECT -4.800 502.940 2.400 504.140 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    PORT
      LAYER met3 ;
        RECT 2917.600 1635.140 2924.800 1636.340 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    PORT
      LAYER met2 ;
        RECT 637.510 3517.600 638.070 3524.800 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    PORT
      LAYER met3 ;
        RECT 2917.600 747.740 2924.800 748.940 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    PORT
      LAYER met2 ;
        RECT 827.490 3517.600 828.050 3524.800 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    PORT
      LAYER met2 ;
        RECT 1191.350 3517.600 1191.910 3524.800 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    PORT
      LAYER met3 ;
        RECT 2917.600 2682.340 2924.800 2683.540 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    PORT
      LAYER met2 ;
        RECT 1716.210 -4.800 1716.770 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    PORT
      LAYER met3 ;
        RECT -4.800 1652.140 2.400 1653.340 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    PORT
      LAYER met2 ;
        RECT 2527.650 3517.600 2528.210 3524.800 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    PORT
      LAYER met2 ;
        RECT 750.210 3517.600 750.770 3524.800 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    PORT
      LAYER met3 ;
        RECT 2917.600 3307.940 2924.800 3309.140 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    PORT
      LAYER met3 ;
        RECT -4.800 3406.540 2.400 3407.740 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    PORT
      LAYER met3 ;
        RECT 2917.600 1835.740 2924.800 1836.940 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    PORT
      LAYER met3 ;
        RECT 2917.600 2240.340 2924.800 2241.540 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    PORT
      LAYER met2 ;
        RECT 476.510 -4.800 477.070 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    PORT
      LAYER met3 ;
        RECT 2917.600 2440.940 2924.800 2442.140 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    PORT
      LAYER met2 ;
        RECT 1258.970 -4.800 1259.530 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    PORT
      LAYER met2 ;
        RECT 1374.890 -4.800 1375.450 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    PORT
      LAYER met3 ;
        RECT -4.800 3022.340 2.400 3023.540 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    PORT
      LAYER met3 ;
        RECT -4.800 2661.940 2.400 2663.140 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    PORT
      LAYER met3 ;
        RECT 2917.600 60.940 2924.800 62.140 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    PORT
      LAYER met3 ;
        RECT -4.800 985.740 2.400 986.940 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    PORT
      LAYER met3 ;
        RECT 2917.600 1573.940 2924.800 1575.140 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    PORT
      LAYER met3 ;
        RECT -4.800 482.540 2.400 483.740 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    PORT
      LAYER met3 ;
        RECT -4.800 2559.940 2.400 2561.140 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    PORT
      LAYER met3 ;
        RECT -4.800 2842.140 2.400 2843.340 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    PORT
      LAYER met2 ;
        RECT 1413.530 -4.800 1414.090 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    PORT
      LAYER met3 ;
        RECT 2917.600 2865.940 2924.800 2867.140 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    PORT
      LAYER met2 ;
        RECT 598.870 3517.600 599.430 3524.800 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    PORT
      LAYER met3 ;
        RECT -4.800 2519.140 2.400 2520.340 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    PORT
      LAYER met2 ;
        RECT 1265.410 3517.600 1265.970 3524.800 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    PORT
      LAYER met2 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    PORT
      LAYER met2 ;
        RECT 846.810 3517.600 847.370 3524.800 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    PORT
      LAYER met3 ;
        RECT 2917.600 1271.340 2924.800 1272.540 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    PORT
      LAYER met2 ;
        RECT 808.170 3517.600 808.730 3524.800 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    PORT
      LAYER met3 ;
        RECT 2917.600 948.340 2924.800 949.540 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    PORT
      LAYER met2 ;
        RECT 763.090 -4.800 763.650 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    PORT
      LAYER met3 ;
        RECT 2917.600 1937.740 2924.800 1938.940 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    PORT
      LAYER met3 ;
        RECT 2917.600 2563.340 2924.800 2564.540 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    PORT
      LAYER met2 ;
        RECT 2546.970 3517.600 2547.530 3524.800 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    PORT
      LAYER met3 ;
        RECT -4.800 1934.340 2.400 1935.540 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    PORT
      LAYER met3 ;
        RECT -4.800 1067.340 2.400 1068.540 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    PORT
      LAYER met3 ;
        RECT -4.800 1410.740 2.400 1411.940 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    PORT
      LAYER met3 ;
        RECT -4.800 3508.540 2.400 3509.740 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    PORT
      LAYER met2 ;
        RECT 1011.030 -4.800 1011.590 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    PORT
      LAYER met2 ;
        RECT 2852.870 3517.600 2853.430 3524.800 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    PORT
      LAYER met2 ;
        RECT 1877.210 3517.600 1877.770 3524.800 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    PORT
      LAYER met2 ;
        RECT 2041.430 -4.800 2041.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    PORT
      LAYER met3 ;
        RECT 2917.600 3226.340 2924.800 3227.540 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    PORT
      LAYER met3 ;
        RECT 2917.600 1958.140 2924.800 1959.340 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    PORT
      LAYER met3 ;
        RECT 2917.600 122.140 2924.800 123.340 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    PORT
      LAYER met2 ;
        RECT 2260.390 3517.600 2260.950 3524.800 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    PORT
      LAYER met2 ;
        RECT 93.330 -4.800 93.890 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    PORT
      LAYER met2 ;
        RECT 924.090 3517.600 924.650 3524.800 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    PORT
      LAYER met2 ;
        RECT 1896.530 3517.600 1897.090 3524.800 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    PORT
      LAYER met3 ;
        RECT -4.800 1148.940 2.400 1150.140 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    PORT
      LAYER met3 ;
        RECT 2917.600 686.540 2924.800 687.740 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    PORT
      LAYER met3 ;
        RECT 2917.600 2400.140 2924.800 2401.340 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    PORT
      LAYER met3 ;
        RECT -4.800 159.540 2.400 160.740 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    PORT
      LAYER met3 ;
        RECT -4.800 1774.540 2.400 1775.740 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    PORT
      LAYER met2 ;
        RECT 1126.950 -4.800 1127.510 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    PORT
      LAYER met3 ;
        RECT 2917.600 203.740 2924.800 204.940 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    PORT
      LAYER met3 ;
        RECT -4.800 1811.940 2.400 1813.140 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    PORT
      LAYER met3 ;
        RECT -4.800 2277.740 2.400 2278.940 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    PORT
      LAYER met2 ;
        RECT 1706.550 3517.600 1707.110 3524.800 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    PORT
      LAYER met3 ;
        RECT 2917.600 2158.740 2924.800 2159.940 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    PORT
      LAYER met2 ;
        RECT 553.790 -4.800 554.350 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    PORT
      LAYER met2 ;
        RECT 940.190 3517.600 940.750 3524.800 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    PORT
      LAYER met3 ;
        RECT 2917.600 465.540 2924.800 466.740 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    PORT
      LAYER met3 ;
        RECT -4.800 139.140 2.400 140.340 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    PORT
      LAYER met3 ;
        RECT 2917.600 1128.540 2924.800 1129.740 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    PORT
      LAYER met3 ;
        RECT 2917.600 3491.540 2924.800 3492.740 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    PORT
      LAYER met3 ;
        RECT 2917.600 1148.940 2924.800 1150.140 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    PORT
      LAYER met3 ;
        RECT -4.800 3447.340 2.400 3448.540 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    PORT
      LAYER met2 ;
        RECT 2347.330 -4.800 2347.890 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    PORT
      LAYER met3 ;
        RECT 2917.600 2338.940 2924.800 2340.140 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    PORT
      LAYER met3 ;
        RECT -4.800 462.140 2.400 463.340 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    PORT
      LAYER met2 ;
        RECT 1545.550 -4.800 1546.110 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    PORT
      LAYER met2 ;
        RECT 1526.230 -4.800 1526.790 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    PORT
      LAYER met2 ;
        RECT 2385.970 -4.800 2386.530 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    PORT
      LAYER met2 ;
        RECT 1362.010 3517.600 1362.570 3524.800 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    PORT
      LAYER met3 ;
        RECT -4.800 1189.740 2.400 1190.940 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    PORT
      LAYER met3 ;
        RECT -4.800 1087.740 2.400 1088.940 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    PORT
      LAYER met3 ;
        RECT 2917.600 1009.540 2924.800 1010.740 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    PORT
      LAYER met2 ;
        RECT 1584.190 -4.800 1584.750 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    PORT
      LAYER met3 ;
        RECT -4.800 1611.340 2.400 1612.540 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    PORT
      LAYER met2 ;
        RECT 2640.350 3517.600 2640.910 3524.800 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    PORT
      LAYER met3 ;
        RECT 2917.600 40.540 2924.800 41.740 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    PORT
      LAYER met3 ;
        RECT 2917.600 343.140 2924.800 344.340 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    PORT
      LAYER met3 ;
        RECT 2917.600 645.740 2924.800 646.940 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    PORT
      LAYER met3 ;
        RECT -4.800 400.940 2.400 402.140 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    PORT
      LAYER met3 ;
        RECT 2917.600 1733.740 2924.800 1734.940 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    PORT
      LAYER met2 ;
        RECT 1857.890 3517.600 1858.450 3524.800 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    PORT
      LAYER met2 ;
        RECT 1226.770 3517.600 1227.330 3524.800 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    PORT
      LAYER met3 ;
        RECT -4.800 3467.740 2.400 3468.940 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    PORT
      LAYER met2 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    PORT
      LAYER met2 ;
        RECT 1890.090 -4.800 1890.650 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    PORT
      LAYER met2 ;
        RECT 424.990 3517.600 425.550 3524.800 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    PORT
      LAYER met3 ;
        RECT -4.800 3144.740 2.400 3145.940 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    PORT
      LAYER met2 ;
        RECT 2807.790 -4.800 2808.350 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    PORT
      LAYER met2 ;
        RECT 730.890 3517.600 731.450 3524.800 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    PORT
      LAYER met2 ;
        RECT 2431.050 3517.600 2431.610 3524.800 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    PORT
      LAYER met3 ;
        RECT -4.800 2155.340 2.400 2156.540 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    PORT
      LAYER met2 ;
        RECT 1851.450 -4.800 1852.010 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    PORT
      LAYER met3 ;
        RECT -4.800 421.340 2.400 422.540 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    PORT
      LAYER met2 ;
        RECT 2202.430 3517.600 2202.990 3524.800 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    PORT
      LAYER met2 ;
        RECT 1986.690 -4.800 1987.250 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    PORT
      LAYER met3 ;
        RECT -4.800 1006.140 2.400 1007.340 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    PORT
      LAYER met2 ;
        RECT 1400.650 3517.600 1401.210 3524.800 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    PORT
      LAYER met2 ;
        RECT 235.010 3517.600 235.570 3524.800 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    PORT
      LAYER met3 ;
        RECT 2917.600 625.340 2924.800 626.540 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    PORT
      LAYER met3 ;
        RECT 2917.600 2138.340 2924.800 2139.540 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    PORT
      LAYER met2 ;
        RECT 1774.170 -4.800 1774.730 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    PORT
      LAYER met3 ;
        RECT -4.800 3226.340 2.400 3227.540 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    PORT
      LAYER met3 ;
        RECT -4.800 2056.740 2.400 2057.940 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    PORT
      LAYER met2 ;
        RECT 1812.810 -4.800 1813.370 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    PORT
      LAYER met2 ;
        RECT 2183.110 3517.600 2183.670 3524.800 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    PORT
      LAYER met3 ;
        RECT -4.800 1369.940 2.400 1371.140 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    PORT
      LAYER met2 ;
        RECT 2614.590 -4.800 2615.150 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    PORT
      LAYER met3 ;
        RECT 2917.600 -0.260 2924.800 0.940 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    PORT
      LAYER met3 ;
        RECT -4.800 744.340 2.400 745.540 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    PORT
      LAYER met3 ;
        RECT -4.800 319.340 2.400 320.540 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    PORT
      LAYER met3 ;
        RECT 2917.600 907.540 2924.800 908.740 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    PORT
      LAYER met2 ;
        RECT 1603.510 -4.800 1604.070 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    PORT
      LAYER met2 ;
        RECT 2366.650 -4.800 2367.210 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    PORT
      LAYER met3 ;
        RECT -4.800 241.140 2.400 242.340 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    PORT
      LAYER met2 ;
        RECT 2221.750 3517.600 2222.310 3524.800 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    PORT
      LAYER met2 ;
        RECT 1793.490 -4.800 1794.050 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    PORT
      LAYER met2 ;
        RECT 25.710 3517.600 26.270 3524.800 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    PORT
      LAYER met2 ;
        RECT 2002.790 -4.800 2003.350 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    PORT
      LAYER met3 ;
        RECT -4.800 3345.340 2.400 3346.540 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    PORT
      LAYER met3 ;
        RECT 2917.600 2379.740 2924.800 2380.940 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    PORT
      LAYER met2 ;
        RECT 1661.470 -4.800 1662.030 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    PORT
      LAYER met3 ;
        RECT 2917.600 768.140 2924.800 769.340 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    PORT
      LAYER met3 ;
        RECT 2917.600 220.740 2924.800 221.940 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    PORT
      LAYER met3 ;
        RECT 2917.600 1169.340 2924.800 1170.540 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    PORT
      LAYER met3 ;
        RECT -4.800 2862.540 2.400 2863.740 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    PORT
      LAYER met2 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    PORT
      LAYER met3 ;
        RECT -4.800 2801.340 2.400 2802.540 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    PORT
      LAYER met2 ;
        RECT 2308.690 -4.800 2309.250 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    PORT
      LAYER met2 ;
        RECT 2585.610 3517.600 2586.170 3524.800 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    PORT
      LAYER met2 ;
        RECT 579.550 3517.600 580.110 3524.800 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    PORT
      LAYER met2 ;
        RECT 2891.510 3517.600 2892.070 3524.800 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    PORT
      LAYER met3 ;
        RECT -4.800 564.140 2.400 565.340 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    PORT
      LAYER met3 ;
        RECT 2917.600 383.940 2924.800 385.140 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    PORT
      LAYER met3 ;
        RECT 2917.600 2199.540 2924.800 2200.740 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    PORT
      LAYER met2 ;
        RECT 1133.390 3517.600 1133.950 3524.800 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    PORT
      LAYER met2 ;
        RECT 2118.710 -4.800 2119.270 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    PORT
      LAYER met2 ;
        RECT 856.470 -4.800 857.030 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    PORT
      LAYER met2 ;
        RECT 2086.510 3517.600 2087.070 3524.800 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    PORT
      LAYER met2 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    PORT
      LAYER met3 ;
        RECT -4.800 1390.340 2.400 1391.540 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    PORT
      LAYER met2 ;
        RECT 45.030 3517.600 45.590 3524.800 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    PORT
      LAYER met2 ;
        RECT 953.070 -4.800 953.630 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    PORT
      LAYER met2 ;
        RECT 2775.590 3517.600 2776.150 3524.800 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    PORT
      LAYER met2 ;
        RECT 2556.630 -4.800 2557.190 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    PORT
      LAYER met3 ;
        RECT 2917.600 1431.140 2924.800 1432.340 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    PORT
      LAYER met2 ;
        RECT 2125.150 3517.600 2125.710 3524.800 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    PORT
      LAYER met3 ;
        RECT -4.800 1046.940 2.400 1048.140 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    PORT
      LAYER met3 ;
        RECT -4.800 2400.140 2.400 2401.340 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    PORT
      LAYER met2 ;
        RECT 1487.590 -4.800 1488.150 2.400 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    PORT
      LAYER met2 ;
        RECT 1754.850 -4.800 1755.410 2.400 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    PORT
      LAYER met2 ;
        RECT 215.690 3517.600 216.250 3524.800 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    PORT
      LAYER met3 ;
        RECT 2917.600 808.940 2924.800 810.140 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    PORT
      LAYER met2 ;
        RECT 2105.830 3517.600 2106.390 3524.800 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    PORT
      LAYER met2 ;
        RECT 840.370 -4.800 840.930 2.400 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    PORT
      LAYER met3 ;
        RECT 2917.600 2359.340 2924.800 2360.540 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    PORT
      LAYER met2 ;
        RECT 885.450 3517.600 886.010 3524.800 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    PORT
      LAYER met2 ;
        RECT 2566.290 3517.600 2566.850 3524.800 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    PORT
      LAYER met2 ;
        RECT 711.570 3517.600 712.130 3524.800 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    PORT
      LAYER met2 ;
        RECT 177.050 3517.600 177.610 3524.800 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    PORT
      LAYER met3 ;
        RECT -4.800 601.540 2.400 602.740 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    PORT
      LAYER met2 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    PORT
      LAYER met3 ;
        RECT 2917.600 2984.940 2924.800 2986.140 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    PORT
      LAYER met2 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    PORT
      LAYER met3 ;
        RECT 2917.600 2179.140 2924.800 2180.340 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    PORT
      LAYER met2 ;
        RECT 627.850 -4.800 628.410 2.400 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    PORT
      LAYER met2 ;
        RECT 1304.050 3517.600 1304.610 3524.800 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    PORT
      LAYER met3 ;
        RECT -4.800 220.740 2.400 221.940 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    PORT
      LAYER met2 ;
        RECT 1700.110 -4.800 1700.670 2.400 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    PORT
      LAYER met2 ;
        RECT 2814.230 3517.600 2814.790 3524.800 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    PORT
      LAYER met3 ;
        RECT -4.800 1893.540 2.400 1894.740 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    PORT
      LAYER met3 ;
        RECT 2917.600 564.140 2924.800 565.340 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    PORT
      LAYER met2 ;
        RECT 64.350 3517.600 64.910 3524.800 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    PORT
      LAYER met2 ;
        RECT 254.330 3517.600 254.890 3524.800 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    PORT
      LAYER met2 ;
        RECT 1181.690 -4.800 1182.250 2.400 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    PORT
      LAYER met2 ;
        RECT 1439.290 3517.600 1439.850 3524.800 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    PORT
      LAYER met3 ;
        RECT 2917.600 3188.940 2924.800 3190.140 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    PORT
      LAYER met3 ;
        RECT 2917.600 1512.740 2924.800 1513.940 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    PORT
      LAYER met3 ;
        RECT -4.800 1590.940 2.400 1592.140 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    PORT
      LAYER met3 ;
        RECT -4.800 965.340 2.400 966.540 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    PORT
      LAYER met3 ;
        RECT 2917.600 1230.540 2924.800 1231.740 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    PORT
      LAYER met3 ;
        RECT -4.800 200.340 2.400 201.540 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    PORT
      LAYER met2 ;
        RECT 1419.970 3517.600 1420.530 3524.800 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    PORT
      LAYER met3 ;
        RECT -4.800 764.740 2.400 765.940 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    PORT
      LAYER met3 ;
        RECT -4.800 360.140 2.400 361.340 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    PORT
      LAYER met2 ;
        RECT 933.750 -4.800 934.310 2.400 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    PORT
      LAYER met3 ;
        RECT 2917.600 968.740 2924.800 969.940 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    PORT
      LAYER met2 ;
        RECT 209.250 -4.800 209.810 2.400 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    PORT
      LAYER met2 ;
        RECT 972.390 -4.800 972.950 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    PORT
      LAYER met3 ;
        RECT 2917.600 887.140 2924.800 888.340 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    PORT
      LAYER met2 ;
        RECT 2910.830 3517.600 2911.390 3524.800 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    PORT
      LAYER met3 ;
        RECT 2917.600 1794.940 2924.800 1796.140 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    PORT
      LAYER met2 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    PORT
      LAYER met3 ;
        RECT 2917.600 1533.140 2924.800 1534.340 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    PORT
      LAYER met3 ;
        RECT -4.800 77.940 2.400 79.140 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    PORT
      LAYER met2 ;
        RECT 2299.030 3517.600 2299.590 3524.800 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    PORT
      LAYER met2 ;
        RECT 2099.390 -4.800 2099.950 2.400 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    PORT
      LAYER met3 ;
        RECT 2917.600 2219.940 2924.800 2221.140 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    PORT
      LAYER met2 ;
        RECT 2698.310 3517.600 2698.870 3524.800 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    PORT
      LAYER met3 ;
        RECT -4.800 118.740 2.400 119.940 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    PORT
      LAYER met2 ;
        RECT 1532.670 3517.600 1533.230 3524.800 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    PORT
      LAYER met2 ;
        RECT 2736.950 3517.600 2737.510 3524.800 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    PORT
      LAYER met2 ;
        RECT 386.350 3517.600 386.910 3524.800 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    PORT
      LAYER met3 ;
        RECT -4.800 1509.340 2.400 1510.540 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    PORT
      LAYER met3 ;
        RECT 2917.600 584.540 2924.800 585.740 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    PORT
      LAYER met3 ;
        RECT -4.800 1451.540 2.400 1452.740 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    PORT
      LAYER met3 ;
        RECT 2917.600 2318.540 2924.800 2319.740 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    PORT
      LAYER met2 ;
        RECT 1075.430 3517.600 1075.990 3524.800 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    PORT
      LAYER met2 ;
        RECT 2501.890 -4.800 2502.450 2.400 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    PORT
      LAYER met3 ;
        RECT 2917.600 3086.940 2924.800 3088.140 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    PORT
      LAYER met3 ;
        RECT 2917.600 2661.940 2924.800 2663.140 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    PORT
      LAYER met2 ;
        RECT 2450.370 3517.600 2450.930 3524.800 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    PORT
      LAYER met3 ;
        RECT 2917.600 3409.940 2924.800 3411.140 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    PORT
      LAYER met3 ;
        RECT 2917.600 81.340 2924.800 82.540 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    PORT
      LAYER met3 ;
        RECT -4.800 57.540 2.400 58.740 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    PORT
      LAYER met2 ;
        RECT 2881.850 -4.800 2882.410 2.400 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    PORT
      LAYER met3 ;
        RECT 2917.600 543.740 2924.800 544.940 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    PORT
      LAYER met2 ;
        RECT 589.210 -4.800 589.770 2.400 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    PORT
      LAYER met2 ;
        RECT 875.790 -4.800 876.350 2.400 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    PORT
      LAYER met3 ;
        RECT 2917.600 183.340 2924.800 184.540 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    PORT
      LAYER met3 ;
        RECT 2917.600 1373.340 2924.800 1374.540 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    PORT
      LAYER met3 ;
        RECT 2917.600 3107.340 2924.800 3108.540 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    PORT
      LAYER met2 ;
        RECT 1172.030 3517.600 1172.590 3524.800 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    PORT
      LAYER met2 ;
        RECT 1017.470 3517.600 1018.030 3524.800 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    PORT
      LAYER met2 ;
        RECT 521.590 3517.600 522.150 3524.800 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    PORT
      LAYER met2 ;
        RECT 1088.310 -4.800 1088.870 2.400 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    PORT
      LAYER met3 ;
        RECT 2917.600 3450.740 2924.800 3451.940 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    PORT
      LAYER met3 ;
        RECT -4.800 904.140 2.400 905.340 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    PORT
      LAYER met2 ;
        RECT 331.610 3517.600 332.170 3524.800 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    PORT
      LAYER met3 ;
        RECT -4.800 261.540 2.400 262.740 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    PORT
      LAYER met3 ;
        RECT 2917.600 3046.140 2924.800 3047.340 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    PORT
      LAYER met2 ;
        RECT 1780.610 3517.600 1781.170 3524.800 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    PORT
      LAYER met2 ;
        RECT 1571.310 3517.600 1571.870 3524.800 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    PORT
      LAYER met2 ;
        RECT 2144.470 3517.600 2145.030 3524.800 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    PORT
      LAYER met2 ;
        RECT 2318.350 3517.600 2318.910 3524.800 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    PORT
      LAYER met2 ;
        RECT 2337.670 3517.600 2338.230 3524.800 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    PORT
      LAYER met3 ;
        RECT -4.800 1206.740 2.400 1207.940 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    PORT
      LAYER met2 ;
        RECT 1246.090 3517.600 1246.650 3524.800 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    PORT
      LAYER met3 ;
        RECT -4.800 1128.540 2.400 1129.740 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    PORT
      LAYER met2 ;
        RECT 35.370 -4.800 35.930 2.400 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    PORT
      LAYER met2 ;
        RECT 2862.530 -4.800 2863.090 2.400 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    PORT
      LAYER met3 ;
        RECT -4.800 1267.940 2.400 1269.140 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    PORT
      LAYER met3 ;
        RECT 2917.600 989.140 2924.800 990.340 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    PORT
      LAYER met3 ;
        RECT -4.800 2216.540 2.400 2217.740 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    PORT
      LAYER met3 ;
        RECT 2917.600 1312.140 2924.800 1313.340 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    PORT
      LAYER met3 ;
        RECT -4.800 2923.740 2.400 2924.940 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    PORT
      LAYER met2 ;
        RECT 151.290 -4.800 151.850 2.400 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    PORT
      LAYER met3 ;
        RECT -4.800 1308.740 2.400 1309.940 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    PORT
      LAYER met3 ;
        RECT -4.800 866.740 2.400 867.940 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    PORT
      LAYER met2 ;
        RECT 1210.670 3517.600 1211.230 3524.800 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    PORT
      LAYER met3 ;
        RECT 2917.600 20.140 2924.800 21.340 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    PORT
      LAYER met2 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    PORT
      LAYER met3 ;
        RECT -4.800 2478.340 2.400 2479.540 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    PORT
      LAYER met3 ;
        RECT 2917.600 2641.540 2924.800 2642.740 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    PORT
      LAYER met3 ;
        RECT 2917.600 3348.740 2924.800 3349.940 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    PORT
      LAYER met2 ;
        RECT 2827.110 -4.800 2827.670 2.400 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    PORT
      LAYER met3 ;
        RECT -4.800 2944.140 2.400 2945.340 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    PORT
      LAYER met3 ;
        RECT 2917.600 706.940 2924.800 708.140 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    PORT
      LAYER met3 ;
        RECT 2917.600 3168.540 2924.800 3169.740 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    PORT
      LAYER met2 ;
        RECT 769.530 3517.600 770.090 3524.800 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    PORT
      LAYER met3 ;
        RECT 2917.600 2702.740 2924.800 2703.940 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    PORT
      LAYER met2 ;
        RECT 2749.830 -4.800 2750.390 2.400 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    PORT
      LAYER met2 ;
        RECT 1551.990 3517.600 1552.550 3524.800 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    PORT
      LAYER met3 ;
        RECT 2917.600 1091.140 2924.800 1092.340 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    PORT
      LAYER met2 ;
        RECT 540.910 3517.600 541.470 3524.800 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    PORT
      LAYER met3 ;
        RECT 2917.600 424.740 2924.800 425.940 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    PORT
      LAYER met3 ;
        RECT -4.800 2114.540 2.400 2115.740 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    PORT
      LAYER met2 ;
        RECT 457.190 -4.800 457.750 2.400 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    PORT
      LAYER met3 ;
        RECT 2917.600 2583.740 2924.800 2584.940 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    PORT
      LAYER met2 ;
        RECT 2022.110 -4.800 2022.670 2.400 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    PORT
      LAYER met3 ;
        RECT -4.800 1108.140 2.400 1109.340 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    PORT
      LAYER met2 ;
        RECT 914.430 -4.800 914.990 2.400 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    PORT
      LAYER met3 ;
        RECT -4.800 1471.940 2.400 1473.140 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    PORT
      LAYER met3 ;
        RECT -4.800 3083.540 2.400 3084.740 ;
    END
  END la_oenb[9]
  PIN user_clock2
    PORT
      LAYER met2 ;
        RECT 1590.630 3517.600 1591.190 3524.800 ;
    END
  END user_clock2
  PIN user_irq[0]
    PORT
      LAYER met3 ;
        RECT 2917.600 3511.940 2924.800 3513.140 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    PORT
      LAYER met3 ;
        RECT -4.800 2984.940 2.400 2986.140 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    PORT
      LAYER met3 ;
        RECT -4.800 3304.540 2.400 3305.740 ;
    END
  END user_irq[2]
  PIN vccd1
    PORT
      LAYER met5 ;
        RECT -43.630 3434.330 2963.250 3437.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3254.330 2963.250 3257.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3074.330 2963.250 3077.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2894.330 2963.250 2897.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2714.330 2963.250 2717.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2534.330 2963.250 2537.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2354.330 2963.250 2357.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2174.330 2963.250 2177.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1994.330 2963.250 1997.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1814.330 2963.250 1817.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1634.330 2963.250 1637.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1454.330 2963.250 1457.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1274.330 2963.250 1277.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1094.330 2963.250 1097.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 914.330 2963.250 917.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 734.330 2963.250 737.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 554.330 2963.250 557.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 374.330 2963.250 377.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 194.330 2963.250 197.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 14.330 2963.250 17.430 ;
    END
    PORT
      LAYER met4 ;
        RECT 2888.970 -38.270 2892.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 -38.270 2712.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 -38.270 2532.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 -38.270 2352.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 -38.270 2172.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1988.970 -38.270 1992.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 -38.270 1812.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1628.970 -38.270 1632.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1448.970 -38.270 1452.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1268.970 -38.270 1272.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.970 -38.270 1092.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.970 -38.270 912.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 -38.270 732.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 -38.270 552.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 -38.270 372.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 -38.270 192.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.970 -38.270 12.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2926.550 -4.670 2929.650 3524.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -10.030 3521.250 2929.650 3524.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -10.030 -4.670 2929.650 -1.570 ;
    END
    PORT
      LAYER met4 ;
        RECT -10.030 -4.670 -6.930 3524.350 ;
    END
  END vccd1
  PIN vccd2
    PORT
      LAYER met5 ;
        RECT -43.630 3471.530 2963.250 3474.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3291.530 2963.250 3294.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3111.530 2963.250 3114.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2931.530 2963.250 2934.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2751.530 2963.250 2754.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2571.530 2963.250 2574.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2391.530 2963.250 2394.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2211.530 2963.250 2214.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2031.530 2963.250 2034.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1851.530 2963.250 1854.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1671.530 2963.250 1674.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1491.530 2963.250 1494.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1311.530 2963.250 1314.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1131.530 2963.250 1134.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 951.530 2963.250 954.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 771.530 2963.250 774.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 591.530 2963.250 594.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 411.530 2963.250 414.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 231.530 2963.250 234.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 51.530 2963.250 54.630 ;
    END
    PORT
      LAYER met4 ;
        RECT 2746.170 -38.270 2749.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2566.170 -38.270 2569.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2386.170 -38.270 2389.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2206.170 -38.270 2209.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2026.170 -38.270 2029.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1846.170 -38.270 1849.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1666.170 -38.270 1669.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1486.170 -38.270 1489.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1306.170 -38.270 1309.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1126.170 -38.270 1129.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 946.170 -38.270 949.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 766.170 -38.270 769.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 586.170 -38.270 589.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 406.170 -38.270 409.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 226.170 -38.270 229.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 46.170 -38.270 49.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2936.150 -14.270 2939.250 3533.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -19.630 3530.850 2939.250 3533.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -19.630 -14.270 2939.250 -11.170 ;
    END
    PORT
      LAYER met4 ;
        RECT -19.630 -14.270 -16.530 3533.950 ;
    END
  END vccd2
  PIN vdda1
    PORT
      LAYER met5 ;
        RECT -43.630 3328.730 2963.250 3331.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3148.730 2963.250 3151.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2968.730 2963.250 2971.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2788.730 2963.250 2791.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2608.730 2963.250 2611.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2428.730 2963.250 2431.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2248.730 2963.250 2251.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2068.730 2963.250 2071.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1888.730 2963.250 1891.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1708.730 2963.250 1711.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1528.730 2963.250 1531.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1348.730 2963.250 1351.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1168.730 2963.250 1171.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 988.730 2963.250 991.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 808.730 2963.250 811.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 628.730 2963.250 631.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 448.730 2963.250 451.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 268.730 2963.250 271.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 88.730 2963.250 91.830 ;
    END
    PORT
      LAYER met4 ;
        RECT 2783.370 -38.270 2786.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2603.370 -38.270 2606.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2423.370 -38.270 2426.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2243.370 -38.270 2246.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2063.370 -38.270 2066.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1883.370 -38.270 1886.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1703.370 -38.270 1706.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1523.370 -38.270 1526.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1343.370 -38.270 1346.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1163.370 -38.270 1166.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 983.370 -38.270 986.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 803.370 -38.270 806.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 623.370 -38.270 626.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 443.370 -38.270 446.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 263.370 -38.270 266.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 83.370 -38.270 86.470 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2945.750 -23.870 2948.850 3543.550 ;
    END
    PORT
      LAYER met5 ;
        RECT -29.230 3540.450 2948.850 3543.550 ;
    END
    PORT
      LAYER met5 ;
        RECT -29.230 -23.870 2948.850 -20.770 ;
    END
    PORT
      LAYER met4 ;
        RECT -29.230 -23.870 -26.130 3543.550 ;
    END
  END vdda1
  PIN vdda2
    PORT
      LAYER met5 ;
        RECT -43.630 3365.930 2963.250 3369.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3185.930 2963.250 3189.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3005.930 2963.250 3009.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2825.930 2963.250 2829.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2645.930 2963.250 2649.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2465.930 2963.250 2469.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2285.930 2963.250 2289.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2105.930 2963.250 2109.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1925.930 2963.250 1929.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1745.930 2963.250 1749.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1565.930 2963.250 1569.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1385.930 2963.250 1389.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1205.930 2963.250 1209.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1025.930 2963.250 1029.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 845.930 2963.250 849.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 665.930 2963.250 669.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 485.930 2963.250 489.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 305.930 2963.250 309.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 125.930 2963.250 129.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 2820.570 -38.270 2823.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2640.570 -38.270 2643.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2460.570 -38.270 2463.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2280.570 -38.270 2283.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2100.570 -38.270 2103.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1920.570 -38.270 1923.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1740.570 -38.270 1743.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1560.570 -38.270 1563.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1380.570 -38.270 1383.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1200.570 -38.270 1203.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1020.570 -38.270 1023.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 840.570 -38.270 843.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 660.570 -38.270 663.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 480.570 -38.270 483.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 300.570 -38.270 303.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 120.570 -38.270 123.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2955.350 -33.470 2958.450 3553.150 ;
    END
    PORT
      LAYER met5 ;
        RECT -38.830 3550.050 2958.450 3553.150 ;
    END
    PORT
      LAYER met5 ;
        RECT -38.830 -33.470 2958.450 -30.370 ;
    END
    PORT
      LAYER met4 ;
        RECT -38.830 -33.470 -35.730 3553.150 ;
    END
  END vdda2
  PIN vssa1
    PORT
      LAYER met5 ;
        RECT -43.630 3347.330 2963.250 3350.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3167.330 2963.250 3170.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2987.330 2963.250 2990.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2807.330 2963.250 2810.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2627.330 2963.250 2630.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2447.330 2963.250 2450.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2267.330 2963.250 2270.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2087.330 2963.250 2090.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1907.330 2963.250 1910.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1727.330 2963.250 1730.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1547.330 2963.250 1550.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1367.330 2963.250 1370.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1187.330 2963.250 1190.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1007.330 2963.250 1010.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 827.330 2963.250 830.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 647.330 2963.250 650.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 467.330 2963.250 470.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 287.330 2963.250 290.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 107.330 2963.250 110.430 ;
    END
    PORT
      LAYER met4 ;
        RECT 2801.970 -38.270 2805.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2621.970 -38.270 2625.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2441.970 -38.270 2445.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2261.970 -38.270 2265.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2081.970 -38.270 2085.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1901.970 -38.270 1905.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1721.970 -38.270 1725.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1541.970 -38.270 1545.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1361.970 -38.270 1365.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1181.970 -38.270 1185.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1001.970 -38.270 1005.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 821.970 -38.270 825.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 641.970 -38.270 645.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 461.970 -38.270 465.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 281.970 -38.270 285.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 101.970 -38.270 105.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2950.550 -28.670 2953.650 3548.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3545.250 2953.650 3548.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 -28.670 2953.650 -25.570 ;
    END
    PORT
      LAYER met4 ;
        RECT -34.030 -28.670 -30.930 3548.350 ;
    END
  END vssa1
  PIN vssa2
    PORT
      LAYER met5 ;
        RECT -43.630 3384.530 2963.250 3387.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3204.530 2963.250 3207.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3024.530 2963.250 3027.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2844.530 2963.250 2847.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2664.530 2963.250 2667.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2484.530 2963.250 2487.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2304.530 2963.250 2307.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2124.530 2963.250 2127.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1944.530 2963.250 1947.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1764.530 2963.250 1767.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1584.530 2963.250 1587.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1404.530 2963.250 1407.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1224.530 2963.250 1227.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1044.530 2963.250 1047.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 864.530 2963.250 867.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 684.530 2963.250 687.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 504.530 2963.250 507.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 324.530 2963.250 327.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 144.530 2963.250 147.630 ;
    END
    PORT
      LAYER met4 ;
        RECT 2839.170 -38.270 2842.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2659.170 -38.270 2662.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2479.170 -38.270 2482.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2299.170 -38.270 2302.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2119.170 -38.270 2122.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1939.170 -38.270 1942.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1759.170 -38.270 1762.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1579.170 -38.270 1582.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1399.170 -38.270 1402.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1219.170 -38.270 1222.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1039.170 -38.270 1042.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 859.170 -38.270 862.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 679.170 -38.270 682.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 499.170 -38.270 502.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 319.170 -38.270 322.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 139.170 -38.270 142.270 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2960.150 -38.270 2963.250 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3554.850 2963.250 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 -38.270 2963.250 -35.170 ;
    END
    PORT
      LAYER met4 ;
        RECT -43.630 -38.270 -40.530 3557.950 ;
    END
  END vssa2
  PIN vssd1
    PORT
      LAYER met5 ;
        RECT -43.630 3452.930 2963.250 3456.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3272.930 2963.250 3276.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3092.930 2963.250 3096.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2912.930 2963.250 2916.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2732.930 2963.250 2736.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2552.930 2963.250 2556.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2372.930 2963.250 2376.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2192.930 2963.250 2196.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2012.930 2963.250 2016.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1832.930 2963.250 1836.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1652.930 2963.250 1656.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1472.930 2963.250 1476.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1292.930 2963.250 1296.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1112.930 2963.250 1116.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 932.930 2963.250 936.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 752.930 2963.250 756.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 572.930 2963.250 576.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 392.930 2963.250 396.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 212.930 2963.250 216.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 32.930 2963.250 36.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 2907.570 -38.270 2910.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2727.570 -38.270 2730.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2547.570 -38.270 2550.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2367.570 -38.270 2370.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2187.570 -38.270 2190.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2007.570 -38.270 2010.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1827.570 -38.270 1830.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1647.570 -38.270 1650.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1467.570 -38.270 1470.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1287.570 -38.270 1290.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1107.570 -38.270 1110.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 927.570 -38.270 930.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 747.570 -38.270 750.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 567.570 -38.270 570.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 387.570 -38.270 390.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 207.570 -38.270 210.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 27.570 -38.270 30.670 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2931.350 -9.470 2934.450 3529.150 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3526.050 2934.450 3529.150 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 -9.470 2934.450 -6.370 ;
    END
    PORT
      LAYER met4 ;
        RECT -14.830 -9.470 -11.730 3529.150 ;
    END
  END vssd1
  PIN vssd2
    PORT
      LAYER met5 ;
        RECT -43.630 3490.130 2963.250 3493.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3310.130 2963.250 3313.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3130.130 2963.250 3133.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2950.130 2963.250 2953.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2770.130 2963.250 2773.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2590.130 2963.250 2593.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2410.130 2963.250 2413.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2230.130 2963.250 2233.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2050.130 2963.250 2053.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1870.130 2963.250 1873.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1690.130 2963.250 1693.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1510.130 2963.250 1513.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1330.130 2963.250 1333.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1150.130 2963.250 1153.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 970.130 2963.250 973.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 790.130 2963.250 793.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 610.130 2963.250 613.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 430.130 2963.250 433.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 250.130 2963.250 253.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 70.130 2963.250 73.230 ;
    END
    PORT
      LAYER met4 ;
        RECT 2764.770 -38.270 2767.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2584.770 -38.270 2587.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2404.770 -38.270 2407.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2224.770 -38.270 2227.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2044.770 -38.270 2047.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.770 -38.270 1867.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1684.770 -38.270 1687.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1504.770 -38.270 1507.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1324.770 -38.270 1327.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1144.770 -38.270 1147.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 964.770 -38.270 967.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 784.770 -38.270 787.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.770 -38.270 607.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 424.770 -38.270 427.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 244.770 -38.270 247.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.770 -38.270 67.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2940.950 -19.070 2944.050 3538.750 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3535.650 2944.050 3538.750 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 -19.070 2944.050 -15.970 ;
    END
    PORT
      LAYER met4 ;
        RECT -24.430 -19.070 -21.330 3538.750 ;
    END
  END vssd2
  PIN wb_clk_i
    PORT
      LAYER met3 ;
        RECT 2917.600 1291.740 2924.800 1292.940 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    PORT
      LAYER met3 ;
        RECT -4.800 1754.140 2.400 1755.340 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    PORT
      LAYER met3 ;
        RECT 2917.600 1917.340 2924.800 1918.540 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    PORT
      LAYER met2 ;
        RECT 998.150 3517.600 998.710 3524.800 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    PORT
      LAYER met2 ;
        RECT 273.650 3517.600 274.210 3524.800 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    PORT
      LAYER met3 ;
        RECT -4.800 2359.340 2.400 2360.540 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    PORT
      LAYER met2 ;
        RECT 321.950 -4.800 322.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    PORT
      LAYER met2 ;
        RECT 1948.050 -4.800 1948.610 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    PORT
      LAYER met3 ;
        RECT 2917.600 3287.540 2924.800 3288.740 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    PORT
      LAYER met3 ;
        RECT 2917.600 3066.540 2924.800 3067.740 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    PORT
      LAYER met2 ;
        RECT 2215.310 -4.800 2215.870 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    PORT
      LAYER met3 ;
        RECT 2917.600 2784.340 2924.800 2785.540 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    PORT
      LAYER met3 ;
        RECT 2917.600 1716.740 2924.800 1717.940 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    PORT
      LAYER met3 ;
        RECT 2917.600 445.140 2924.800 446.340 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    PORT
      LAYER met2 ;
        RECT 1036.790 3517.600 1037.350 3524.800 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    PORT
      LAYER met2 ;
        RECT 2031.770 3517.600 2032.330 3524.800 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    PORT
      LAYER met2 ;
        RECT 1967.370 -4.800 1967.930 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    PORT
      LAYER met2 ;
        RECT 2788.470 -4.800 2789.030 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    PORT
      LAYER met3 ;
        RECT 2917.600 1393.740 2924.800 1394.940 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    PORT
      LAYER met3 ;
        RECT -4.800 2780.940 2.400 2782.140 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    PORT
      LAYER met2 ;
        RECT 1870.770 -4.800 1871.330 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    PORT
      LAYER met2 ;
        RECT 360.590 -4.800 361.150 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    PORT
      LAYER met3 ;
        RECT -4.800 98.340 2.400 99.540 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    PORT
      LAYER met3 ;
        RECT 2917.600 2621.140 2924.800 2622.340 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    PORT
      LAYER met2 ;
        RECT 2489.010 3517.600 2489.570 3524.800 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    PORT
      LAYER met2 ;
        RECT 1336.250 -4.800 1336.810 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    PORT
      LAYER met2 ;
        RECT 1667.910 3517.600 1668.470 3524.800 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    PORT
      LAYER met3 ;
        RECT 2917.600 2019.340 2924.800 2020.540 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    PORT
      LAYER met2 ;
        RECT 2653.230 -4.800 2653.790 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    PORT
      LAYER met2 ;
        RECT 1609.950 3517.600 1610.510 3524.800 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    PORT
      LAYER met3 ;
        RECT -4.800 543.740 2.400 544.940 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    PORT
      LAYER met2 ;
        RECT 1068.990 -4.800 1069.550 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    PORT
      LAYER met2 ;
        RECT 170.610 -4.800 171.170 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    PORT
      LAYER met3 ;
        RECT 2917.600 485.940 2924.800 487.140 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    PORT
      LAYER met3 ;
        RECT 2917.600 1451.540 2924.800 1452.740 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    PORT
      LAYER met2 ;
        RECT 157.730 3517.600 158.290 3524.800 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    PORT
      LAYER met2 ;
        RECT 2872.190 3517.600 2872.750 3524.800 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    PORT
      LAYER met3 ;
        RECT -4.800 1794.940 2.400 1796.140 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    PORT
      LAYER met3 ;
        RECT -4.800 2036.340 2.400 2037.540 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    PORT
      LAYER met3 ;
        RECT -4.800 1954.740 2.400 1955.940 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    PORT
      LAYER met2 ;
        RECT 131.970 -4.800 132.530 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    PORT
      LAYER met2 ;
        RECT 724.450 -4.800 725.010 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    PORT
      LAYER met3 ;
        RECT 2917.600 2281.140 2924.800 2282.340 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    PORT
      LAYER met2 ;
        RECT 1928.730 -4.800 1929.290 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    PORT
      LAYER met2 ;
        RECT 1458.610 3517.600 1459.170 3524.800 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    PORT
      LAYER met2 ;
        RECT 2279.710 3517.600 2280.270 3524.800 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    PORT
      LAYER met3 ;
        RECT -4.800 2882.940 2.400 2884.140 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    PORT
      LAYER met2 ;
        RECT 515.150 -4.800 515.710 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    PORT
      LAYER met3 ;
        RECT 2917.600 2542.940 2924.800 2544.140 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    PORT
      LAYER met2 ;
        RECT 2411.730 3517.600 2412.290 3524.800 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    PORT
      LAYER met3 ;
        RECT -4.800 1329.140 2.400 1330.340 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    PORT
      LAYER met3 ;
        RECT 2917.600 3148.140 2924.800 3149.340 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    PORT
      LAYER met3 ;
        RECT 2917.600 1553.540 2924.800 1554.740 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    PORT
      LAYER met2 ;
        RECT 2289.370 -4.800 2289.930 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    PORT
      LAYER met2 ;
        RECT 2051.090 3517.600 2051.650 3524.800 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    PORT
      LAYER met2 ;
        RECT 99.770 3517.600 100.330 3524.800 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    PORT
      LAYER met2 ;
        RECT 1030.350 -4.800 1030.910 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    PORT
      LAYER met3 ;
        RECT 2917.600 2481.740 2924.800 2482.940 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    PORT
      LAYER met2 ;
        RECT 2691.870 -4.800 2692.430 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    PORT
      LAYER met3 ;
        RECT 2917.600 1414.140 2924.800 1415.340 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    PORT
      LAYER met3 ;
        RECT -4.800 1247.540 2.400 1248.740 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    PORT
      LAYER met3 ;
        RECT 2917.600 506.340 2924.800 507.540 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    PORT
      LAYER met2 ;
        RECT 534.470 -4.800 535.030 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    PORT
      LAYER met2 ;
        RECT 1622.830 -4.800 1623.390 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    PORT
      LAYER met3 ;
        RECT -4.800 16.740 2.400 17.940 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    PORT
      LAYER met2 ;
        RECT 1993.130 3517.600 1993.690 3524.800 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    PORT
      LAYER met3 ;
        RECT 2917.600 3430.340 2924.800 3431.540 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    PORT
      LAYER met3 ;
        RECT 2917.600 523.340 2924.800 524.540 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    PORT
      LAYER met2 ;
        RECT 267.210 -4.800 267.770 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    PORT
      LAYER met3 ;
        RECT 2917.600 2301.540 2924.800 2302.740 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    PORT
      LAYER met2 ;
        RECT 74.010 -4.800 74.570 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    PORT
      LAYER met3 ;
        RECT 2917.600 3471.140 2924.800 3472.340 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    PORT
      LAYER met2 ;
        RECT 1915.850 3517.600 1916.410 3524.800 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    PORT
      LAYER met3 ;
        RECT 2917.600 727.340 2924.800 728.540 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    PORT
      LAYER met2 ;
        RECT 1819.250 3517.600 1819.810 3524.800 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    PORT
      LAYER met3 ;
        RECT -4.800 584.540 2.400 585.740 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    PORT
      LAYER met3 ;
        RECT -4.800 683.140 2.400 684.340 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    PORT
      LAYER met2 ;
        RECT 2176.670 -4.800 2177.230 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    PORT
      LAYER met2 ;
        RECT -0.050 -4.800 0.510 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    PORT
      LAYER met2 ;
        RECT 2540.530 -4.800 2541.090 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    PORT
      LAYER met3 ;
        RECT -4.800 1288.340 2.400 1289.540 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    PORT
      LAYER met3 ;
        RECT -4.800 2621.140 2.400 2622.340 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    PORT
      LAYER met2 ;
        RECT 463.630 3517.600 464.190 3524.800 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    PORT
      LAYER met3 ;
        RECT -4.800 846.340 2.400 847.540 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    PORT
      LAYER met2 ;
        RECT 666.490 -4.800 667.050 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    PORT
      LAYER met2 ;
        RECT 247.890 -4.800 248.450 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    PORT
      LAYER met2 ;
        RECT 1284.730 3517.600 1285.290 3524.800 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    PORT
      LAYER met2 ;
        RECT 560.230 3517.600 560.790 3524.800 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    PORT
      LAYER met2 ;
        RECT 1735.530 -4.800 1736.090 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    PORT
      LAYER met2 ;
        RECT 1838.570 3517.600 1839.130 3524.800 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    PORT
      LAYER met3 ;
        RECT 2917.600 1210.140 2924.800 1211.340 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    PORT
      LAYER met3 ;
        RECT -4.800 2015.940 2.400 2017.140 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    PORT
      LAYER met3 ;
        RECT 2917.600 2845.540 2924.800 2846.740 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    PORT
      LAYER met2 ;
        RECT 705.130 -4.800 705.690 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    PORT
      LAYER met2 ;
        RECT 1220.330 -4.800 1220.890 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    PORT
      LAYER met3 ;
        RECT -4.800 179.940 2.400 181.140 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    PORT
      LAYER met3 ;
        RECT 2917.600 2723.140 2924.800 2724.340 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    PORT
      LAYER met2 ;
        RECT 1909.410 -4.800 1909.970 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    PORT
      LAYER met2 ;
        RECT 1799.930 3517.600 1800.490 3524.800 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    PORT
      LAYER met2 ;
        RECT 1764.510 3517.600 1765.070 3524.800 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    PORT
      LAYER met3 ;
        RECT -4.800 3001.940 2.400 3003.140 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    PORT
      LAYER met2 ;
        RECT 80.450 3517.600 81.010 3524.800 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    PORT
      LAYER met2 ;
        RECT 2273.270 -4.800 2273.830 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    PORT
      LAYER met3 ;
        RECT -4.800 703.540 2.400 704.740 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    PORT
      LAYER met3 ;
        RECT -4.800 2719.740 2.400 2720.940 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    PORT
      LAYER met3 ;
        RECT 2917.600 1856.140 2924.800 1857.340 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2914.100 3508.885 ;
      LAYER met1 ;
        RECT 2.830 6.840 2914.950 3511.480 ;
      LAYER met2 ;
        RECT 0.090 3517.320 6.110 3518.050 ;
        RECT 7.230 3517.320 25.430 3518.050 ;
        RECT 26.550 3517.320 44.750 3518.050 ;
        RECT 45.870 3517.320 64.070 3518.050 ;
        RECT 65.190 3517.320 80.170 3518.050 ;
        RECT 81.290 3517.320 99.490 3518.050 ;
        RECT 100.610 3517.320 118.810 3518.050 ;
        RECT 119.930 3517.320 138.130 3518.050 ;
        RECT 139.250 3517.320 157.450 3518.050 ;
        RECT 158.570 3517.320 176.770 3518.050 ;
        RECT 177.890 3517.320 196.090 3518.050 ;
        RECT 197.210 3517.320 215.410 3518.050 ;
        RECT 216.530 3517.320 234.730 3518.050 ;
        RECT 235.850 3517.320 254.050 3518.050 ;
        RECT 255.170 3517.320 273.370 3518.050 ;
        RECT 274.490 3517.320 292.690 3518.050 ;
        RECT 293.810 3517.320 312.010 3518.050 ;
        RECT 313.130 3517.320 331.330 3518.050 ;
        RECT 332.450 3517.320 350.650 3518.050 ;
        RECT 351.770 3517.320 366.750 3518.050 ;
        RECT 367.870 3517.320 386.070 3518.050 ;
        RECT 387.190 3517.320 405.390 3518.050 ;
        RECT 406.510 3517.320 424.710 3518.050 ;
        RECT 425.830 3517.320 444.030 3518.050 ;
        RECT 445.150 3517.320 463.350 3518.050 ;
        RECT 464.470 3517.320 482.670 3518.050 ;
        RECT 483.790 3517.320 501.990 3518.050 ;
        RECT 503.110 3517.320 521.310 3518.050 ;
        RECT 522.430 3517.320 540.630 3518.050 ;
        RECT 541.750 3517.320 559.950 3518.050 ;
        RECT 561.070 3517.320 579.270 3518.050 ;
        RECT 580.390 3517.320 598.590 3518.050 ;
        RECT 599.710 3517.320 617.910 3518.050 ;
        RECT 619.030 3517.320 637.230 3518.050 ;
        RECT 638.350 3517.320 653.330 3518.050 ;
        RECT 654.450 3517.320 672.650 3518.050 ;
        RECT 673.770 3517.320 691.970 3518.050 ;
        RECT 693.090 3517.320 711.290 3518.050 ;
        RECT 712.410 3517.320 730.610 3518.050 ;
        RECT 731.730 3517.320 749.930 3518.050 ;
        RECT 751.050 3517.320 769.250 3518.050 ;
        RECT 770.370 3517.320 788.570 3518.050 ;
        RECT 789.690 3517.320 807.890 3518.050 ;
        RECT 809.010 3517.320 827.210 3518.050 ;
        RECT 828.330 3517.320 846.530 3518.050 ;
        RECT 847.650 3517.320 865.850 3518.050 ;
        RECT 866.970 3517.320 885.170 3518.050 ;
        RECT 886.290 3517.320 904.490 3518.050 ;
        RECT 905.610 3517.320 923.810 3518.050 ;
        RECT 924.930 3517.320 939.910 3518.050 ;
        RECT 941.030 3517.320 959.230 3518.050 ;
        RECT 960.350 3517.320 978.550 3518.050 ;
        RECT 979.670 3517.320 997.870 3518.050 ;
        RECT 998.990 3517.320 1017.190 3518.050 ;
        RECT 1018.310 3517.320 1036.510 3518.050 ;
        RECT 1037.630 3517.320 1055.830 3518.050 ;
        RECT 1056.950 3517.320 1075.150 3518.050 ;
        RECT 1076.270 3517.320 1094.470 3518.050 ;
        RECT 1095.590 3517.320 1113.790 3518.050 ;
        RECT 1114.910 3517.320 1133.110 3518.050 ;
        RECT 1134.230 3517.320 1152.430 3518.050 ;
        RECT 1153.550 3517.320 1171.750 3518.050 ;
        RECT 1172.870 3517.320 1191.070 3518.050 ;
        RECT 1192.190 3517.320 1210.390 3518.050 ;
        RECT 1211.510 3517.320 1226.490 3518.050 ;
        RECT 1227.610 3517.320 1245.810 3518.050 ;
        RECT 1246.930 3517.320 1265.130 3518.050 ;
        RECT 1266.250 3517.320 1284.450 3518.050 ;
        RECT 1285.570 3517.320 1303.770 3518.050 ;
        RECT 1304.890 3517.320 1323.090 3518.050 ;
        RECT 1324.210 3517.320 1342.410 3518.050 ;
        RECT 1343.530 3517.320 1361.730 3518.050 ;
        RECT 1362.850 3517.320 1381.050 3518.050 ;
        RECT 1382.170 3517.320 1400.370 3518.050 ;
        RECT 1401.490 3517.320 1419.690 3518.050 ;
        RECT 1420.810 3517.320 1439.010 3518.050 ;
        RECT 1440.130 3517.320 1458.330 3518.050 ;
        RECT 1459.450 3517.320 1477.650 3518.050 ;
        RECT 1478.770 3517.320 1496.970 3518.050 ;
        RECT 1498.090 3517.320 1513.070 3518.050 ;
        RECT 1514.190 3517.320 1532.390 3518.050 ;
        RECT 1533.510 3517.320 1551.710 3518.050 ;
        RECT 1552.830 3517.320 1571.030 3518.050 ;
        RECT 1572.150 3517.320 1590.350 3518.050 ;
        RECT 1591.470 3517.320 1609.670 3518.050 ;
        RECT 1610.790 3517.320 1628.990 3518.050 ;
        RECT 1630.110 3517.320 1648.310 3518.050 ;
        RECT 1649.430 3517.320 1667.630 3518.050 ;
        RECT 1668.750 3517.320 1686.950 3518.050 ;
        RECT 1688.070 3517.320 1706.270 3518.050 ;
        RECT 1707.390 3517.320 1725.590 3518.050 ;
        RECT 1726.710 3517.320 1744.910 3518.050 ;
        RECT 1746.030 3517.320 1764.230 3518.050 ;
        RECT 1765.350 3517.320 1780.330 3518.050 ;
        RECT 1781.450 3517.320 1799.650 3518.050 ;
        RECT 1800.770 3517.320 1818.970 3518.050 ;
        RECT 1820.090 3517.320 1838.290 3518.050 ;
        RECT 1839.410 3517.320 1857.610 3518.050 ;
        RECT 1858.730 3517.320 1876.930 3518.050 ;
        RECT 1878.050 3517.320 1896.250 3518.050 ;
        RECT 1897.370 3517.320 1915.570 3518.050 ;
        RECT 1916.690 3517.320 1934.890 3518.050 ;
        RECT 1936.010 3517.320 1954.210 3518.050 ;
        RECT 1955.330 3517.320 1973.530 3518.050 ;
        RECT 1974.650 3517.320 1992.850 3518.050 ;
        RECT 1993.970 3517.320 2012.170 3518.050 ;
        RECT 2013.290 3517.320 2031.490 3518.050 ;
        RECT 2032.610 3517.320 2050.810 3518.050 ;
        RECT 2051.930 3517.320 2066.910 3518.050 ;
        RECT 2068.030 3517.320 2086.230 3518.050 ;
        RECT 2087.350 3517.320 2105.550 3518.050 ;
        RECT 2106.670 3517.320 2124.870 3518.050 ;
        RECT 2125.990 3517.320 2144.190 3518.050 ;
        RECT 2145.310 3517.320 2163.510 3518.050 ;
        RECT 2164.630 3517.320 2182.830 3518.050 ;
        RECT 2183.950 3517.320 2202.150 3518.050 ;
        RECT 2203.270 3517.320 2221.470 3518.050 ;
        RECT 2222.590 3517.320 2240.790 3518.050 ;
        RECT 2241.910 3517.320 2260.110 3518.050 ;
        RECT 2261.230 3517.320 2279.430 3518.050 ;
        RECT 2280.550 3517.320 2298.750 3518.050 ;
        RECT 2299.870 3517.320 2318.070 3518.050 ;
        RECT 2319.190 3517.320 2337.390 3518.050 ;
        RECT 2338.510 3517.320 2353.490 3518.050 ;
        RECT 2354.610 3517.320 2372.810 3518.050 ;
        RECT 2373.930 3517.320 2392.130 3518.050 ;
        RECT 2393.250 3517.320 2411.450 3518.050 ;
        RECT 2412.570 3517.320 2430.770 3518.050 ;
        RECT 2431.890 3517.320 2450.090 3518.050 ;
        RECT 2451.210 3517.320 2469.410 3518.050 ;
        RECT 2470.530 3517.320 2488.730 3518.050 ;
        RECT 2489.850 3517.320 2508.050 3518.050 ;
        RECT 2509.170 3517.320 2527.370 3518.050 ;
        RECT 2528.490 3517.320 2546.690 3518.050 ;
        RECT 2547.810 3517.320 2566.010 3518.050 ;
        RECT 2567.130 3517.320 2585.330 3518.050 ;
        RECT 2586.450 3517.320 2604.650 3518.050 ;
        RECT 2605.770 3517.320 2623.970 3518.050 ;
        RECT 2625.090 3517.320 2640.070 3518.050 ;
        RECT 2641.190 3517.320 2659.390 3518.050 ;
        RECT 2660.510 3517.320 2678.710 3518.050 ;
        RECT 2679.830 3517.320 2698.030 3518.050 ;
        RECT 2699.150 3517.320 2717.350 3518.050 ;
        RECT 2718.470 3517.320 2736.670 3518.050 ;
        RECT 2737.790 3517.320 2755.990 3518.050 ;
        RECT 2757.110 3517.320 2775.310 3518.050 ;
        RECT 2776.430 3517.320 2794.630 3518.050 ;
        RECT 2795.750 3517.320 2813.950 3518.050 ;
        RECT 2815.070 3517.320 2833.270 3518.050 ;
        RECT 2834.390 3517.320 2852.590 3518.050 ;
        RECT 2853.710 3517.320 2871.910 3518.050 ;
        RECT 2873.030 3517.320 2891.230 3518.050 ;
        RECT 2892.350 3517.320 2910.550 3518.050 ;
        RECT 2911.670 3517.320 2914.920 3518.050 ;
        RECT 0.090 2.680 2914.920 3517.320 ;
        RECT 0.790 0.155 15.770 2.680 ;
        RECT 16.890 0.155 35.090 2.680 ;
        RECT 36.210 0.155 54.410 2.680 ;
        RECT 55.530 0.155 73.730 2.680 ;
        RECT 74.850 0.155 93.050 2.680 ;
        RECT 94.170 0.155 112.370 2.680 ;
        RECT 113.490 0.155 131.690 2.680 ;
        RECT 132.810 0.155 151.010 2.680 ;
        RECT 152.130 0.155 170.330 2.680 ;
        RECT 171.450 0.155 189.650 2.680 ;
        RECT 190.770 0.155 208.970 2.680 ;
        RECT 210.090 0.155 228.290 2.680 ;
        RECT 229.410 0.155 247.610 2.680 ;
        RECT 248.730 0.155 266.930 2.680 ;
        RECT 268.050 0.155 283.030 2.680 ;
        RECT 284.150 0.155 302.350 2.680 ;
        RECT 303.470 0.155 321.670 2.680 ;
        RECT 322.790 0.155 340.990 2.680 ;
        RECT 342.110 0.155 360.310 2.680 ;
        RECT 361.430 0.155 379.630 2.680 ;
        RECT 380.750 0.155 398.950 2.680 ;
        RECT 400.070 0.155 418.270 2.680 ;
        RECT 419.390 0.155 437.590 2.680 ;
        RECT 438.710 0.155 456.910 2.680 ;
        RECT 458.030 0.155 476.230 2.680 ;
        RECT 477.350 0.155 495.550 2.680 ;
        RECT 496.670 0.155 514.870 2.680 ;
        RECT 515.990 0.155 534.190 2.680 ;
        RECT 535.310 0.155 553.510 2.680 ;
        RECT 554.630 0.155 569.610 2.680 ;
        RECT 570.730 0.155 588.930 2.680 ;
        RECT 590.050 0.155 608.250 2.680 ;
        RECT 609.370 0.155 627.570 2.680 ;
        RECT 628.690 0.155 646.890 2.680 ;
        RECT 648.010 0.155 666.210 2.680 ;
        RECT 667.330 0.155 685.530 2.680 ;
        RECT 686.650 0.155 704.850 2.680 ;
        RECT 705.970 0.155 724.170 2.680 ;
        RECT 725.290 0.155 743.490 2.680 ;
        RECT 744.610 0.155 762.810 2.680 ;
        RECT 763.930 0.155 782.130 2.680 ;
        RECT 783.250 0.155 801.450 2.680 ;
        RECT 802.570 0.155 820.770 2.680 ;
        RECT 821.890 0.155 840.090 2.680 ;
        RECT 841.210 0.155 856.190 2.680 ;
        RECT 857.310 0.155 875.510 2.680 ;
        RECT 876.630 0.155 894.830 2.680 ;
        RECT 895.950 0.155 914.150 2.680 ;
        RECT 915.270 0.155 933.470 2.680 ;
        RECT 934.590 0.155 952.790 2.680 ;
        RECT 953.910 0.155 972.110 2.680 ;
        RECT 973.230 0.155 991.430 2.680 ;
        RECT 992.550 0.155 1010.750 2.680 ;
        RECT 1011.870 0.155 1030.070 2.680 ;
        RECT 1031.190 0.155 1049.390 2.680 ;
        RECT 1050.510 0.155 1068.710 2.680 ;
        RECT 1069.830 0.155 1088.030 2.680 ;
        RECT 1089.150 0.155 1107.350 2.680 ;
        RECT 1108.470 0.155 1126.670 2.680 ;
        RECT 1127.790 0.155 1142.770 2.680 ;
        RECT 1143.890 0.155 1162.090 2.680 ;
        RECT 1163.210 0.155 1181.410 2.680 ;
        RECT 1182.530 0.155 1200.730 2.680 ;
        RECT 1201.850 0.155 1220.050 2.680 ;
        RECT 1221.170 0.155 1239.370 2.680 ;
        RECT 1240.490 0.155 1258.690 2.680 ;
        RECT 1259.810 0.155 1278.010 2.680 ;
        RECT 1279.130 0.155 1297.330 2.680 ;
        RECT 1298.450 0.155 1316.650 2.680 ;
        RECT 1317.770 0.155 1335.970 2.680 ;
        RECT 1337.090 0.155 1355.290 2.680 ;
        RECT 1356.410 0.155 1374.610 2.680 ;
        RECT 1375.730 0.155 1393.930 2.680 ;
        RECT 1395.050 0.155 1413.250 2.680 ;
        RECT 1414.370 0.155 1429.350 2.680 ;
        RECT 1430.470 0.155 1448.670 2.680 ;
        RECT 1449.790 0.155 1467.990 2.680 ;
        RECT 1469.110 0.155 1487.310 2.680 ;
        RECT 1488.430 0.155 1506.630 2.680 ;
        RECT 1507.750 0.155 1525.950 2.680 ;
        RECT 1527.070 0.155 1545.270 2.680 ;
        RECT 1546.390 0.155 1564.590 2.680 ;
        RECT 1565.710 0.155 1583.910 2.680 ;
        RECT 1585.030 0.155 1603.230 2.680 ;
        RECT 1604.350 0.155 1622.550 2.680 ;
        RECT 1623.670 0.155 1641.870 2.680 ;
        RECT 1642.990 0.155 1661.190 2.680 ;
        RECT 1662.310 0.155 1680.510 2.680 ;
        RECT 1681.630 0.155 1699.830 2.680 ;
        RECT 1700.950 0.155 1715.930 2.680 ;
        RECT 1717.050 0.155 1735.250 2.680 ;
        RECT 1736.370 0.155 1754.570 2.680 ;
        RECT 1755.690 0.155 1773.890 2.680 ;
        RECT 1775.010 0.155 1793.210 2.680 ;
        RECT 1794.330 0.155 1812.530 2.680 ;
        RECT 1813.650 0.155 1831.850 2.680 ;
        RECT 1832.970 0.155 1851.170 2.680 ;
        RECT 1852.290 0.155 1870.490 2.680 ;
        RECT 1871.610 0.155 1889.810 2.680 ;
        RECT 1890.930 0.155 1909.130 2.680 ;
        RECT 1910.250 0.155 1928.450 2.680 ;
        RECT 1929.570 0.155 1947.770 2.680 ;
        RECT 1948.890 0.155 1967.090 2.680 ;
        RECT 1968.210 0.155 1986.410 2.680 ;
        RECT 1987.530 0.155 2002.510 2.680 ;
        RECT 2003.630 0.155 2021.830 2.680 ;
        RECT 2022.950 0.155 2041.150 2.680 ;
        RECT 2042.270 0.155 2060.470 2.680 ;
        RECT 2061.590 0.155 2079.790 2.680 ;
        RECT 2080.910 0.155 2099.110 2.680 ;
        RECT 2100.230 0.155 2118.430 2.680 ;
        RECT 2119.550 0.155 2137.750 2.680 ;
        RECT 2138.870 0.155 2157.070 2.680 ;
        RECT 2158.190 0.155 2176.390 2.680 ;
        RECT 2177.510 0.155 2195.710 2.680 ;
        RECT 2196.830 0.155 2215.030 2.680 ;
        RECT 2216.150 0.155 2234.350 2.680 ;
        RECT 2235.470 0.155 2253.670 2.680 ;
        RECT 2254.790 0.155 2272.990 2.680 ;
        RECT 2274.110 0.155 2289.090 2.680 ;
        RECT 2290.210 0.155 2308.410 2.680 ;
        RECT 2309.530 0.155 2327.730 2.680 ;
        RECT 2328.850 0.155 2347.050 2.680 ;
        RECT 2348.170 0.155 2366.370 2.680 ;
        RECT 2367.490 0.155 2385.690 2.680 ;
        RECT 2386.810 0.155 2405.010 2.680 ;
        RECT 2406.130 0.155 2424.330 2.680 ;
        RECT 2425.450 0.155 2443.650 2.680 ;
        RECT 2444.770 0.155 2462.970 2.680 ;
        RECT 2464.090 0.155 2482.290 2.680 ;
        RECT 2483.410 0.155 2501.610 2.680 ;
        RECT 2502.730 0.155 2520.930 2.680 ;
        RECT 2522.050 0.155 2540.250 2.680 ;
        RECT 2541.370 0.155 2556.350 2.680 ;
        RECT 2557.470 0.155 2575.670 2.680 ;
        RECT 2576.790 0.155 2594.990 2.680 ;
        RECT 2596.110 0.155 2614.310 2.680 ;
        RECT 2615.430 0.155 2633.630 2.680 ;
        RECT 2634.750 0.155 2652.950 2.680 ;
        RECT 2654.070 0.155 2672.270 2.680 ;
        RECT 2673.390 0.155 2691.590 2.680 ;
        RECT 2692.710 0.155 2710.910 2.680 ;
        RECT 2712.030 0.155 2730.230 2.680 ;
        RECT 2731.350 0.155 2749.550 2.680 ;
        RECT 2750.670 0.155 2768.870 2.680 ;
        RECT 2769.990 0.155 2788.190 2.680 ;
        RECT 2789.310 0.155 2807.510 2.680 ;
        RECT 2808.630 0.155 2826.830 2.680 ;
        RECT 2827.950 0.155 2842.930 2.680 ;
        RECT 2844.050 0.155 2862.250 2.680 ;
        RECT 2863.370 0.155 2881.570 2.680 ;
        RECT 2882.690 0.155 2900.890 2.680 ;
        RECT 2902.010 0.155 2914.920 2.680 ;
      LAYER met3 ;
        RECT 0.065 3511.540 2917.200 3512.705 ;
        RECT 0.065 3510.140 2917.930 3511.540 ;
        RECT 2.800 3508.140 2917.930 3510.140 ;
        RECT 0.065 3493.140 2917.930 3508.140 ;
        RECT 0.065 3491.140 2917.200 3493.140 ;
        RECT 0.065 3489.740 2917.930 3491.140 ;
        RECT 2.800 3487.740 2917.930 3489.740 ;
        RECT 0.065 3472.740 2917.930 3487.740 ;
        RECT 0.065 3470.740 2917.200 3472.740 ;
        RECT 0.065 3469.340 2917.930 3470.740 ;
        RECT 2.800 3467.340 2917.930 3469.340 ;
        RECT 0.065 3452.340 2917.930 3467.340 ;
        RECT 0.065 3450.340 2917.200 3452.340 ;
        RECT 0.065 3448.940 2917.930 3450.340 ;
        RECT 2.800 3446.940 2917.930 3448.940 ;
        RECT 0.065 3431.940 2917.930 3446.940 ;
        RECT 0.065 3429.940 2917.200 3431.940 ;
        RECT 0.065 3428.540 2917.930 3429.940 ;
        RECT 2.800 3426.540 2917.930 3428.540 ;
        RECT 0.065 3411.540 2917.930 3426.540 ;
        RECT 0.065 3409.540 2917.200 3411.540 ;
        RECT 0.065 3408.140 2917.930 3409.540 ;
        RECT 2.800 3406.140 2917.930 3408.140 ;
        RECT 0.065 3391.140 2917.930 3406.140 ;
        RECT 0.065 3389.140 2917.200 3391.140 ;
        RECT 0.065 3387.740 2917.930 3389.140 ;
        RECT 2.800 3385.740 2917.930 3387.740 ;
        RECT 0.065 3370.740 2917.930 3385.740 ;
        RECT 0.065 3368.740 2917.200 3370.740 ;
        RECT 0.065 3367.340 2917.930 3368.740 ;
        RECT 2.800 3365.340 2917.930 3367.340 ;
        RECT 0.065 3350.340 2917.930 3365.340 ;
        RECT 0.065 3348.340 2917.200 3350.340 ;
        RECT 0.065 3346.940 2917.930 3348.340 ;
        RECT 2.800 3344.940 2917.930 3346.940 ;
        RECT 0.065 3329.940 2917.930 3344.940 ;
        RECT 0.065 3327.940 2917.200 3329.940 ;
        RECT 0.065 3326.540 2917.930 3327.940 ;
        RECT 2.800 3324.540 2917.930 3326.540 ;
        RECT 0.065 3309.540 2917.930 3324.540 ;
        RECT 0.065 3307.540 2917.200 3309.540 ;
        RECT 0.065 3306.140 2917.930 3307.540 ;
        RECT 2.800 3304.140 2917.930 3306.140 ;
        RECT 0.065 3289.140 2917.930 3304.140 ;
        RECT 2.800 3287.140 2917.200 3289.140 ;
        RECT 0.065 3268.740 2917.930 3287.140 ;
        RECT 2.800 3266.740 2917.200 3268.740 ;
        RECT 0.065 3248.340 2917.930 3266.740 ;
        RECT 2.800 3246.340 2917.200 3248.340 ;
        RECT 0.065 3227.940 2917.930 3246.340 ;
        RECT 2.800 3225.940 2917.200 3227.940 ;
        RECT 0.065 3210.940 2917.930 3225.940 ;
        RECT 0.065 3208.940 2917.200 3210.940 ;
        RECT 0.065 3207.540 2917.930 3208.940 ;
        RECT 2.800 3205.540 2917.930 3207.540 ;
        RECT 0.065 3190.540 2917.930 3205.540 ;
        RECT 0.065 3188.540 2917.200 3190.540 ;
        RECT 0.065 3187.140 2917.930 3188.540 ;
        RECT 2.800 3185.140 2917.930 3187.140 ;
        RECT 0.065 3170.140 2917.930 3185.140 ;
        RECT 0.065 3168.140 2917.200 3170.140 ;
        RECT 0.065 3166.740 2917.930 3168.140 ;
        RECT 2.800 3164.740 2917.930 3166.740 ;
        RECT 0.065 3149.740 2917.930 3164.740 ;
        RECT 0.065 3147.740 2917.200 3149.740 ;
        RECT 0.065 3146.340 2917.930 3147.740 ;
        RECT 2.800 3144.340 2917.930 3146.340 ;
        RECT 0.065 3129.340 2917.930 3144.340 ;
        RECT 0.065 3127.340 2917.200 3129.340 ;
        RECT 0.065 3125.940 2917.930 3127.340 ;
        RECT 2.800 3123.940 2917.930 3125.940 ;
        RECT 0.065 3108.940 2917.930 3123.940 ;
        RECT 0.065 3106.940 2917.200 3108.940 ;
        RECT 0.065 3105.540 2917.930 3106.940 ;
        RECT 2.800 3103.540 2917.930 3105.540 ;
        RECT 0.065 3088.540 2917.930 3103.540 ;
        RECT 0.065 3086.540 2917.200 3088.540 ;
        RECT 0.065 3085.140 2917.930 3086.540 ;
        RECT 2.800 3083.140 2917.930 3085.140 ;
        RECT 0.065 3068.140 2917.930 3083.140 ;
        RECT 0.065 3066.140 2917.200 3068.140 ;
        RECT 0.065 3064.740 2917.930 3066.140 ;
        RECT 2.800 3062.740 2917.930 3064.740 ;
        RECT 0.065 3047.740 2917.930 3062.740 ;
        RECT 0.065 3045.740 2917.200 3047.740 ;
        RECT 0.065 3044.340 2917.930 3045.740 ;
        RECT 2.800 3042.340 2917.930 3044.340 ;
        RECT 0.065 3027.340 2917.930 3042.340 ;
        RECT 0.065 3025.340 2917.200 3027.340 ;
        RECT 0.065 3023.940 2917.930 3025.340 ;
        RECT 2.800 3021.940 2917.930 3023.940 ;
        RECT 0.065 3006.940 2917.930 3021.940 ;
        RECT 0.065 3004.940 2917.200 3006.940 ;
        RECT 0.065 3003.540 2917.930 3004.940 ;
        RECT 2.800 3001.540 2917.930 3003.540 ;
        RECT 0.065 2986.540 2917.930 3001.540 ;
        RECT 2.800 2984.540 2917.200 2986.540 ;
        RECT 0.065 2966.140 2917.930 2984.540 ;
        RECT 2.800 2964.140 2917.200 2966.140 ;
        RECT 0.065 2945.740 2917.930 2964.140 ;
        RECT 2.800 2943.740 2917.200 2945.740 ;
        RECT 0.065 2925.340 2917.930 2943.740 ;
        RECT 2.800 2923.340 2917.200 2925.340 ;
        RECT 0.065 2908.340 2917.930 2923.340 ;
        RECT 0.065 2906.340 2917.200 2908.340 ;
        RECT 0.065 2904.940 2917.930 2906.340 ;
        RECT 2.800 2902.940 2917.930 2904.940 ;
        RECT 0.065 2887.940 2917.930 2902.940 ;
        RECT 0.065 2885.940 2917.200 2887.940 ;
        RECT 0.065 2884.540 2917.930 2885.940 ;
        RECT 2.800 2882.540 2917.930 2884.540 ;
        RECT 0.065 2867.540 2917.930 2882.540 ;
        RECT 0.065 2865.540 2917.200 2867.540 ;
        RECT 0.065 2864.140 2917.930 2865.540 ;
        RECT 2.800 2862.140 2917.930 2864.140 ;
        RECT 0.065 2847.140 2917.930 2862.140 ;
        RECT 0.065 2845.140 2917.200 2847.140 ;
        RECT 0.065 2843.740 2917.930 2845.140 ;
        RECT 2.800 2841.740 2917.930 2843.740 ;
        RECT 0.065 2826.740 2917.930 2841.740 ;
        RECT 0.065 2824.740 2917.200 2826.740 ;
        RECT 0.065 2823.340 2917.930 2824.740 ;
        RECT 2.800 2821.340 2917.930 2823.340 ;
        RECT 0.065 2806.340 2917.930 2821.340 ;
        RECT 0.065 2804.340 2917.200 2806.340 ;
        RECT 0.065 2802.940 2917.930 2804.340 ;
        RECT 2.800 2800.940 2917.930 2802.940 ;
        RECT 0.065 2785.940 2917.930 2800.940 ;
        RECT 0.065 2783.940 2917.200 2785.940 ;
        RECT 0.065 2782.540 2917.930 2783.940 ;
        RECT 2.800 2780.540 2917.930 2782.540 ;
        RECT 0.065 2765.540 2917.930 2780.540 ;
        RECT 0.065 2763.540 2917.200 2765.540 ;
        RECT 0.065 2762.140 2917.930 2763.540 ;
        RECT 2.800 2760.140 2917.930 2762.140 ;
        RECT 0.065 2745.140 2917.930 2760.140 ;
        RECT 0.065 2743.140 2917.200 2745.140 ;
        RECT 0.065 2741.740 2917.930 2743.140 ;
        RECT 2.800 2739.740 2917.930 2741.740 ;
        RECT 0.065 2724.740 2917.930 2739.740 ;
        RECT 0.065 2722.740 2917.200 2724.740 ;
        RECT 0.065 2721.340 2917.930 2722.740 ;
        RECT 2.800 2719.340 2917.930 2721.340 ;
        RECT 0.065 2704.340 2917.930 2719.340 ;
        RECT 0.065 2702.340 2917.200 2704.340 ;
        RECT 0.065 2700.940 2917.930 2702.340 ;
        RECT 2.800 2698.940 2917.930 2700.940 ;
        RECT 0.065 2683.940 2917.930 2698.940 ;
        RECT 2.800 2681.940 2917.200 2683.940 ;
        RECT 0.065 2663.540 2917.930 2681.940 ;
        RECT 2.800 2661.540 2917.200 2663.540 ;
        RECT 0.065 2643.140 2917.930 2661.540 ;
        RECT 2.800 2641.140 2917.200 2643.140 ;
        RECT 0.065 2622.740 2917.930 2641.140 ;
        RECT 2.800 2620.740 2917.200 2622.740 ;
        RECT 0.065 2605.740 2917.930 2620.740 ;
        RECT 0.065 2603.740 2917.200 2605.740 ;
        RECT 0.065 2602.340 2917.930 2603.740 ;
        RECT 2.800 2600.340 2917.930 2602.340 ;
        RECT 0.065 2585.340 2917.930 2600.340 ;
        RECT 0.065 2583.340 2917.200 2585.340 ;
        RECT 0.065 2581.940 2917.930 2583.340 ;
        RECT 2.800 2579.940 2917.930 2581.940 ;
        RECT 0.065 2564.940 2917.930 2579.940 ;
        RECT 0.065 2562.940 2917.200 2564.940 ;
        RECT 0.065 2561.540 2917.930 2562.940 ;
        RECT 2.800 2559.540 2917.930 2561.540 ;
        RECT 0.065 2544.540 2917.930 2559.540 ;
        RECT 0.065 2542.540 2917.200 2544.540 ;
        RECT 0.065 2541.140 2917.930 2542.540 ;
        RECT 2.800 2539.140 2917.930 2541.140 ;
        RECT 0.065 2524.140 2917.930 2539.140 ;
        RECT 0.065 2522.140 2917.200 2524.140 ;
        RECT 0.065 2520.740 2917.930 2522.140 ;
        RECT 2.800 2518.740 2917.930 2520.740 ;
        RECT 0.065 2503.740 2917.930 2518.740 ;
        RECT 0.065 2501.740 2917.200 2503.740 ;
        RECT 0.065 2500.340 2917.930 2501.740 ;
        RECT 2.800 2498.340 2917.930 2500.340 ;
        RECT 0.065 2483.340 2917.930 2498.340 ;
        RECT 0.065 2481.340 2917.200 2483.340 ;
        RECT 0.065 2479.940 2917.930 2481.340 ;
        RECT 2.800 2477.940 2917.930 2479.940 ;
        RECT 0.065 2462.940 2917.930 2477.940 ;
        RECT 0.065 2460.940 2917.200 2462.940 ;
        RECT 0.065 2459.540 2917.930 2460.940 ;
        RECT 2.800 2457.540 2917.930 2459.540 ;
        RECT 0.065 2442.540 2917.930 2457.540 ;
        RECT 0.065 2440.540 2917.200 2442.540 ;
        RECT 0.065 2439.140 2917.930 2440.540 ;
        RECT 2.800 2437.140 2917.930 2439.140 ;
        RECT 0.065 2422.140 2917.930 2437.140 ;
        RECT 0.065 2420.140 2917.200 2422.140 ;
        RECT 0.065 2418.740 2917.930 2420.140 ;
        RECT 2.800 2416.740 2917.930 2418.740 ;
        RECT 0.065 2401.740 2917.930 2416.740 ;
        RECT 2.800 2399.740 2917.200 2401.740 ;
        RECT 0.065 2381.340 2917.930 2399.740 ;
        RECT 2.800 2379.340 2917.200 2381.340 ;
        RECT 0.065 2360.940 2917.930 2379.340 ;
        RECT 2.800 2358.940 2917.200 2360.940 ;
        RECT 0.065 2340.540 2917.930 2358.940 ;
        RECT 2.800 2338.540 2917.200 2340.540 ;
        RECT 0.065 2320.140 2917.930 2338.540 ;
        RECT 2.800 2318.140 2917.200 2320.140 ;
        RECT 0.065 2303.140 2917.930 2318.140 ;
        RECT 0.065 2301.140 2917.200 2303.140 ;
        RECT 0.065 2299.740 2917.930 2301.140 ;
        RECT 2.800 2297.740 2917.930 2299.740 ;
        RECT 0.065 2282.740 2917.930 2297.740 ;
        RECT 0.065 2280.740 2917.200 2282.740 ;
        RECT 0.065 2279.340 2917.930 2280.740 ;
        RECT 2.800 2277.340 2917.930 2279.340 ;
        RECT 0.065 2262.340 2917.930 2277.340 ;
        RECT 0.065 2260.340 2917.200 2262.340 ;
        RECT 0.065 2258.940 2917.930 2260.340 ;
        RECT 2.800 2256.940 2917.930 2258.940 ;
        RECT 0.065 2241.940 2917.930 2256.940 ;
        RECT 0.065 2239.940 2917.200 2241.940 ;
        RECT 0.065 2238.540 2917.930 2239.940 ;
        RECT 2.800 2236.540 2917.930 2238.540 ;
        RECT 0.065 2221.540 2917.930 2236.540 ;
        RECT 0.065 2219.540 2917.200 2221.540 ;
        RECT 0.065 2218.140 2917.930 2219.540 ;
        RECT 2.800 2216.140 2917.930 2218.140 ;
        RECT 0.065 2201.140 2917.930 2216.140 ;
        RECT 0.065 2199.140 2917.200 2201.140 ;
        RECT 0.065 2197.740 2917.930 2199.140 ;
        RECT 2.800 2195.740 2917.930 2197.740 ;
        RECT 0.065 2180.740 2917.930 2195.740 ;
        RECT 0.065 2178.740 2917.200 2180.740 ;
        RECT 0.065 2177.340 2917.930 2178.740 ;
        RECT 2.800 2175.340 2917.930 2177.340 ;
        RECT 0.065 2160.340 2917.930 2175.340 ;
        RECT 0.065 2158.340 2917.200 2160.340 ;
        RECT 0.065 2156.940 2917.930 2158.340 ;
        RECT 2.800 2154.940 2917.930 2156.940 ;
        RECT 0.065 2139.940 2917.930 2154.940 ;
        RECT 0.065 2137.940 2917.200 2139.940 ;
        RECT 0.065 2136.540 2917.930 2137.940 ;
        RECT 2.800 2134.540 2917.930 2136.540 ;
        RECT 0.065 2119.540 2917.930 2134.540 ;
        RECT 0.065 2117.540 2917.200 2119.540 ;
        RECT 0.065 2116.140 2917.930 2117.540 ;
        RECT 2.800 2114.140 2917.930 2116.140 ;
        RECT 0.065 2099.140 2917.930 2114.140 ;
        RECT 2.800 2097.140 2917.200 2099.140 ;
        RECT 0.065 2078.740 2917.930 2097.140 ;
        RECT 2.800 2076.740 2917.200 2078.740 ;
        RECT 0.065 2058.340 2917.930 2076.740 ;
        RECT 2.800 2056.340 2917.200 2058.340 ;
        RECT 0.065 2037.940 2917.930 2056.340 ;
        RECT 2.800 2035.940 2917.200 2037.940 ;
        RECT 0.065 2020.940 2917.930 2035.940 ;
        RECT 0.065 2018.940 2917.200 2020.940 ;
        RECT 0.065 2017.540 2917.930 2018.940 ;
        RECT 2.800 2015.540 2917.930 2017.540 ;
        RECT 0.065 2000.540 2917.930 2015.540 ;
        RECT 0.065 1998.540 2917.200 2000.540 ;
        RECT 0.065 1997.140 2917.930 1998.540 ;
        RECT 2.800 1995.140 2917.930 1997.140 ;
        RECT 0.065 1980.140 2917.930 1995.140 ;
        RECT 0.065 1978.140 2917.200 1980.140 ;
        RECT 0.065 1976.740 2917.930 1978.140 ;
        RECT 2.800 1974.740 2917.930 1976.740 ;
        RECT 0.065 1959.740 2917.930 1974.740 ;
        RECT 0.065 1957.740 2917.200 1959.740 ;
        RECT 0.065 1956.340 2917.930 1957.740 ;
        RECT 2.800 1954.340 2917.930 1956.340 ;
        RECT 0.065 1939.340 2917.930 1954.340 ;
        RECT 0.065 1937.340 2917.200 1939.340 ;
        RECT 0.065 1935.940 2917.930 1937.340 ;
        RECT 2.800 1933.940 2917.930 1935.940 ;
        RECT 0.065 1918.940 2917.930 1933.940 ;
        RECT 0.065 1916.940 2917.200 1918.940 ;
        RECT 0.065 1915.540 2917.930 1916.940 ;
        RECT 2.800 1913.540 2917.930 1915.540 ;
        RECT 0.065 1898.540 2917.930 1913.540 ;
        RECT 0.065 1896.540 2917.200 1898.540 ;
        RECT 0.065 1895.140 2917.930 1896.540 ;
        RECT 2.800 1893.140 2917.930 1895.140 ;
        RECT 0.065 1878.140 2917.930 1893.140 ;
        RECT 0.065 1876.140 2917.200 1878.140 ;
        RECT 0.065 1874.740 2917.930 1876.140 ;
        RECT 2.800 1872.740 2917.930 1874.740 ;
        RECT 0.065 1857.740 2917.930 1872.740 ;
        RECT 0.065 1855.740 2917.200 1857.740 ;
        RECT 0.065 1854.340 2917.930 1855.740 ;
        RECT 2.800 1852.340 2917.930 1854.340 ;
        RECT 0.065 1837.340 2917.930 1852.340 ;
        RECT 0.065 1835.340 2917.200 1837.340 ;
        RECT 0.065 1833.940 2917.930 1835.340 ;
        RECT 2.800 1831.940 2917.930 1833.940 ;
        RECT 0.065 1816.940 2917.930 1831.940 ;
        RECT 0.065 1814.940 2917.200 1816.940 ;
        RECT 0.065 1813.540 2917.930 1814.940 ;
        RECT 2.800 1811.540 2917.930 1813.540 ;
        RECT 0.065 1796.540 2917.930 1811.540 ;
        RECT 2.800 1794.540 2917.200 1796.540 ;
        RECT 0.065 1776.140 2917.930 1794.540 ;
        RECT 2.800 1774.140 2917.200 1776.140 ;
        RECT 0.065 1755.740 2917.930 1774.140 ;
        RECT 2.800 1753.740 2917.200 1755.740 ;
        RECT 0.065 1735.340 2917.930 1753.740 ;
        RECT 2.800 1733.340 2917.200 1735.340 ;
        RECT 0.065 1718.340 2917.930 1733.340 ;
        RECT 0.065 1716.340 2917.200 1718.340 ;
        RECT 0.065 1714.940 2917.930 1716.340 ;
        RECT 2.800 1712.940 2917.930 1714.940 ;
        RECT 0.065 1697.940 2917.930 1712.940 ;
        RECT 0.065 1695.940 2917.200 1697.940 ;
        RECT 0.065 1694.540 2917.930 1695.940 ;
        RECT 2.800 1692.540 2917.930 1694.540 ;
        RECT 0.065 1677.540 2917.930 1692.540 ;
        RECT 0.065 1675.540 2917.200 1677.540 ;
        RECT 0.065 1674.140 2917.930 1675.540 ;
        RECT 2.800 1672.140 2917.930 1674.140 ;
        RECT 0.065 1657.140 2917.930 1672.140 ;
        RECT 0.065 1655.140 2917.200 1657.140 ;
        RECT 0.065 1653.740 2917.930 1655.140 ;
        RECT 2.800 1651.740 2917.930 1653.740 ;
        RECT 0.065 1636.740 2917.930 1651.740 ;
        RECT 0.065 1634.740 2917.200 1636.740 ;
        RECT 0.065 1633.340 2917.930 1634.740 ;
        RECT 2.800 1631.340 2917.930 1633.340 ;
        RECT 0.065 1616.340 2917.930 1631.340 ;
        RECT 0.065 1614.340 2917.200 1616.340 ;
        RECT 0.065 1612.940 2917.930 1614.340 ;
        RECT 2.800 1610.940 2917.930 1612.940 ;
        RECT 0.065 1595.940 2917.930 1610.940 ;
        RECT 0.065 1593.940 2917.200 1595.940 ;
        RECT 0.065 1592.540 2917.930 1593.940 ;
        RECT 2.800 1590.540 2917.930 1592.540 ;
        RECT 0.065 1575.540 2917.930 1590.540 ;
        RECT 0.065 1573.540 2917.200 1575.540 ;
        RECT 0.065 1572.140 2917.930 1573.540 ;
        RECT 2.800 1570.140 2917.930 1572.140 ;
        RECT 0.065 1555.140 2917.930 1570.140 ;
        RECT 0.065 1553.140 2917.200 1555.140 ;
        RECT 0.065 1551.740 2917.930 1553.140 ;
        RECT 2.800 1549.740 2917.930 1551.740 ;
        RECT 0.065 1534.740 2917.930 1549.740 ;
        RECT 0.065 1532.740 2917.200 1534.740 ;
        RECT 0.065 1531.340 2917.930 1532.740 ;
        RECT 2.800 1529.340 2917.930 1531.340 ;
        RECT 0.065 1514.340 2917.930 1529.340 ;
        RECT 0.065 1512.340 2917.200 1514.340 ;
        RECT 0.065 1510.940 2917.930 1512.340 ;
        RECT 2.800 1508.940 2917.930 1510.940 ;
        RECT 0.065 1493.940 2917.930 1508.940 ;
        RECT 2.800 1491.940 2917.200 1493.940 ;
        RECT 0.065 1473.540 2917.930 1491.940 ;
        RECT 2.800 1471.540 2917.200 1473.540 ;
        RECT 0.065 1453.140 2917.930 1471.540 ;
        RECT 2.800 1451.140 2917.200 1453.140 ;
        RECT 0.065 1432.740 2917.930 1451.140 ;
        RECT 2.800 1430.740 2917.200 1432.740 ;
        RECT 0.065 1415.740 2917.930 1430.740 ;
        RECT 0.065 1413.740 2917.200 1415.740 ;
        RECT 0.065 1412.340 2917.930 1413.740 ;
        RECT 2.800 1410.340 2917.930 1412.340 ;
        RECT 0.065 1395.340 2917.930 1410.340 ;
        RECT 0.065 1393.340 2917.200 1395.340 ;
        RECT 0.065 1391.940 2917.930 1393.340 ;
        RECT 2.800 1389.940 2917.930 1391.940 ;
        RECT 0.065 1374.940 2917.930 1389.940 ;
        RECT 0.065 1372.940 2917.200 1374.940 ;
        RECT 0.065 1371.540 2917.930 1372.940 ;
        RECT 2.800 1369.540 2917.930 1371.540 ;
        RECT 0.065 1354.540 2917.930 1369.540 ;
        RECT 0.065 1352.540 2917.200 1354.540 ;
        RECT 0.065 1351.140 2917.930 1352.540 ;
        RECT 2.800 1349.140 2917.930 1351.140 ;
        RECT 0.065 1334.140 2917.930 1349.140 ;
        RECT 0.065 1332.140 2917.200 1334.140 ;
        RECT 0.065 1330.740 2917.930 1332.140 ;
        RECT 2.800 1328.740 2917.930 1330.740 ;
        RECT 0.065 1313.740 2917.930 1328.740 ;
        RECT 0.065 1311.740 2917.200 1313.740 ;
        RECT 0.065 1310.340 2917.930 1311.740 ;
        RECT 2.800 1308.340 2917.930 1310.340 ;
        RECT 0.065 1293.340 2917.930 1308.340 ;
        RECT 0.065 1291.340 2917.200 1293.340 ;
        RECT 0.065 1289.940 2917.930 1291.340 ;
        RECT 2.800 1287.940 2917.930 1289.940 ;
        RECT 0.065 1272.940 2917.930 1287.940 ;
        RECT 0.065 1270.940 2917.200 1272.940 ;
        RECT 0.065 1269.540 2917.930 1270.940 ;
        RECT 2.800 1267.540 2917.930 1269.540 ;
        RECT 0.065 1252.540 2917.930 1267.540 ;
        RECT 0.065 1250.540 2917.200 1252.540 ;
        RECT 0.065 1249.140 2917.930 1250.540 ;
        RECT 2.800 1247.140 2917.930 1249.140 ;
        RECT 0.065 1232.140 2917.930 1247.140 ;
        RECT 0.065 1230.140 2917.200 1232.140 ;
        RECT 0.065 1228.740 2917.930 1230.140 ;
        RECT 2.800 1226.740 2917.930 1228.740 ;
        RECT 0.065 1211.740 2917.930 1226.740 ;
        RECT 0.065 1209.740 2917.200 1211.740 ;
        RECT 0.065 1208.340 2917.930 1209.740 ;
        RECT 2.800 1206.340 2917.930 1208.340 ;
        RECT 0.065 1191.340 2917.930 1206.340 ;
        RECT 2.800 1189.340 2917.200 1191.340 ;
        RECT 0.065 1170.940 2917.930 1189.340 ;
        RECT 2.800 1168.940 2917.200 1170.940 ;
        RECT 0.065 1150.540 2917.930 1168.940 ;
        RECT 2.800 1148.540 2917.200 1150.540 ;
        RECT 0.065 1130.140 2917.930 1148.540 ;
        RECT 2.800 1128.140 2917.200 1130.140 ;
        RECT 0.065 1113.140 2917.930 1128.140 ;
        RECT 0.065 1111.140 2917.200 1113.140 ;
        RECT 0.065 1109.740 2917.930 1111.140 ;
        RECT 2.800 1107.740 2917.930 1109.740 ;
        RECT 0.065 1092.740 2917.930 1107.740 ;
        RECT 0.065 1090.740 2917.200 1092.740 ;
        RECT 0.065 1089.340 2917.930 1090.740 ;
        RECT 2.800 1087.340 2917.930 1089.340 ;
        RECT 0.065 1072.340 2917.930 1087.340 ;
        RECT 0.065 1070.340 2917.200 1072.340 ;
        RECT 0.065 1068.940 2917.930 1070.340 ;
        RECT 2.800 1066.940 2917.930 1068.940 ;
        RECT 0.065 1051.940 2917.930 1066.940 ;
        RECT 0.065 1049.940 2917.200 1051.940 ;
        RECT 0.065 1048.540 2917.930 1049.940 ;
        RECT 2.800 1046.540 2917.930 1048.540 ;
        RECT 0.065 1031.540 2917.930 1046.540 ;
        RECT 0.065 1029.540 2917.200 1031.540 ;
        RECT 0.065 1028.140 2917.930 1029.540 ;
        RECT 2.800 1026.140 2917.930 1028.140 ;
        RECT 0.065 1011.140 2917.930 1026.140 ;
        RECT 0.065 1009.140 2917.200 1011.140 ;
        RECT 0.065 1007.740 2917.930 1009.140 ;
        RECT 2.800 1005.740 2917.930 1007.740 ;
        RECT 0.065 990.740 2917.930 1005.740 ;
        RECT 0.065 988.740 2917.200 990.740 ;
        RECT 0.065 987.340 2917.930 988.740 ;
        RECT 2.800 985.340 2917.930 987.340 ;
        RECT 0.065 970.340 2917.930 985.340 ;
        RECT 0.065 968.340 2917.200 970.340 ;
        RECT 0.065 966.940 2917.930 968.340 ;
        RECT 2.800 964.940 2917.930 966.940 ;
        RECT 0.065 949.940 2917.930 964.940 ;
        RECT 0.065 947.940 2917.200 949.940 ;
        RECT 0.065 946.540 2917.930 947.940 ;
        RECT 2.800 944.540 2917.930 946.540 ;
        RECT 0.065 929.540 2917.930 944.540 ;
        RECT 0.065 927.540 2917.200 929.540 ;
        RECT 0.065 926.140 2917.930 927.540 ;
        RECT 2.800 924.140 2917.930 926.140 ;
        RECT 0.065 909.140 2917.930 924.140 ;
        RECT 0.065 907.140 2917.200 909.140 ;
        RECT 0.065 905.740 2917.930 907.140 ;
        RECT 2.800 903.740 2917.930 905.740 ;
        RECT 0.065 888.740 2917.930 903.740 ;
        RECT 2.800 886.740 2917.200 888.740 ;
        RECT 0.065 868.340 2917.930 886.740 ;
        RECT 2.800 866.340 2917.200 868.340 ;
        RECT 0.065 847.940 2917.930 866.340 ;
        RECT 2.800 845.940 2917.200 847.940 ;
        RECT 0.065 827.540 2917.930 845.940 ;
        RECT 2.800 825.540 2917.200 827.540 ;
        RECT 0.065 810.540 2917.930 825.540 ;
        RECT 0.065 808.540 2917.200 810.540 ;
        RECT 0.065 807.140 2917.930 808.540 ;
        RECT 2.800 805.140 2917.930 807.140 ;
        RECT 0.065 790.140 2917.930 805.140 ;
        RECT 0.065 788.140 2917.200 790.140 ;
        RECT 0.065 786.740 2917.930 788.140 ;
        RECT 2.800 784.740 2917.930 786.740 ;
        RECT 0.065 769.740 2917.930 784.740 ;
        RECT 0.065 767.740 2917.200 769.740 ;
        RECT 0.065 766.340 2917.930 767.740 ;
        RECT 2.800 764.340 2917.930 766.340 ;
        RECT 0.065 749.340 2917.930 764.340 ;
        RECT 0.065 747.340 2917.200 749.340 ;
        RECT 0.065 745.940 2917.930 747.340 ;
        RECT 2.800 743.940 2917.930 745.940 ;
        RECT 0.065 728.940 2917.930 743.940 ;
        RECT 0.065 726.940 2917.200 728.940 ;
        RECT 0.065 725.540 2917.930 726.940 ;
        RECT 2.800 723.540 2917.930 725.540 ;
        RECT 0.065 708.540 2917.930 723.540 ;
        RECT 0.065 706.540 2917.200 708.540 ;
        RECT 0.065 705.140 2917.930 706.540 ;
        RECT 2.800 703.140 2917.930 705.140 ;
        RECT 0.065 688.140 2917.930 703.140 ;
        RECT 0.065 686.140 2917.200 688.140 ;
        RECT 0.065 684.740 2917.930 686.140 ;
        RECT 2.800 682.740 2917.930 684.740 ;
        RECT 0.065 667.740 2917.930 682.740 ;
        RECT 0.065 665.740 2917.200 667.740 ;
        RECT 0.065 664.340 2917.930 665.740 ;
        RECT 2.800 662.340 2917.930 664.340 ;
        RECT 0.065 647.340 2917.930 662.340 ;
        RECT 0.065 645.340 2917.200 647.340 ;
        RECT 0.065 643.940 2917.930 645.340 ;
        RECT 2.800 641.940 2917.930 643.940 ;
        RECT 0.065 626.940 2917.930 641.940 ;
        RECT 0.065 624.940 2917.200 626.940 ;
        RECT 0.065 623.540 2917.930 624.940 ;
        RECT 2.800 621.540 2917.930 623.540 ;
        RECT 0.065 606.540 2917.930 621.540 ;
        RECT 0.065 604.540 2917.200 606.540 ;
        RECT 0.065 603.140 2917.930 604.540 ;
        RECT 2.800 601.140 2917.930 603.140 ;
        RECT 0.065 586.140 2917.930 601.140 ;
        RECT 2.800 584.140 2917.200 586.140 ;
        RECT 0.065 565.740 2917.930 584.140 ;
        RECT 2.800 563.740 2917.200 565.740 ;
        RECT 0.065 545.340 2917.930 563.740 ;
        RECT 2.800 543.340 2917.200 545.340 ;
        RECT 0.065 524.940 2917.930 543.340 ;
        RECT 2.800 522.940 2917.200 524.940 ;
        RECT 0.065 507.940 2917.930 522.940 ;
        RECT 0.065 505.940 2917.200 507.940 ;
        RECT 0.065 504.540 2917.930 505.940 ;
        RECT 2.800 502.540 2917.930 504.540 ;
        RECT 0.065 487.540 2917.930 502.540 ;
        RECT 0.065 485.540 2917.200 487.540 ;
        RECT 0.065 484.140 2917.930 485.540 ;
        RECT 2.800 482.140 2917.930 484.140 ;
        RECT 0.065 467.140 2917.930 482.140 ;
        RECT 0.065 465.140 2917.200 467.140 ;
        RECT 0.065 463.740 2917.930 465.140 ;
        RECT 2.800 461.740 2917.930 463.740 ;
        RECT 0.065 446.740 2917.930 461.740 ;
        RECT 0.065 444.740 2917.200 446.740 ;
        RECT 0.065 443.340 2917.930 444.740 ;
        RECT 2.800 441.340 2917.930 443.340 ;
        RECT 0.065 426.340 2917.930 441.340 ;
        RECT 0.065 424.340 2917.200 426.340 ;
        RECT 0.065 422.940 2917.930 424.340 ;
        RECT 2.800 420.940 2917.930 422.940 ;
        RECT 0.065 405.940 2917.930 420.940 ;
        RECT 0.065 403.940 2917.200 405.940 ;
        RECT 0.065 402.540 2917.930 403.940 ;
        RECT 2.800 400.540 2917.930 402.540 ;
        RECT 0.065 385.540 2917.930 400.540 ;
        RECT 0.065 383.540 2917.200 385.540 ;
        RECT 0.065 382.140 2917.930 383.540 ;
        RECT 2.800 380.140 2917.930 382.140 ;
        RECT 0.065 365.140 2917.930 380.140 ;
        RECT 0.065 363.140 2917.200 365.140 ;
        RECT 0.065 361.740 2917.930 363.140 ;
        RECT 2.800 359.740 2917.930 361.740 ;
        RECT 0.065 344.740 2917.930 359.740 ;
        RECT 0.065 342.740 2917.200 344.740 ;
        RECT 0.065 341.340 2917.930 342.740 ;
        RECT 2.800 339.340 2917.930 341.340 ;
        RECT 0.065 324.340 2917.930 339.340 ;
        RECT 0.065 322.340 2917.200 324.340 ;
        RECT 0.065 320.940 2917.930 322.340 ;
        RECT 2.800 318.940 2917.930 320.940 ;
        RECT 0.065 303.940 2917.930 318.940 ;
        RECT 0.065 301.940 2917.200 303.940 ;
        RECT 0.065 300.540 2917.930 301.940 ;
        RECT 2.800 298.540 2917.930 300.540 ;
        RECT 0.065 283.540 2917.930 298.540 ;
        RECT 2.800 281.540 2917.200 283.540 ;
        RECT 0.065 263.140 2917.930 281.540 ;
        RECT 2.800 261.140 2917.200 263.140 ;
        RECT 0.065 242.740 2917.930 261.140 ;
        RECT 2.800 240.740 2917.200 242.740 ;
        RECT 0.065 222.340 2917.930 240.740 ;
        RECT 2.800 220.340 2917.200 222.340 ;
        RECT 0.065 205.340 2917.930 220.340 ;
        RECT 0.065 203.340 2917.200 205.340 ;
        RECT 0.065 201.940 2917.930 203.340 ;
        RECT 2.800 199.940 2917.930 201.940 ;
        RECT 0.065 184.940 2917.930 199.940 ;
        RECT 0.065 182.940 2917.200 184.940 ;
        RECT 0.065 181.540 2917.930 182.940 ;
        RECT 2.800 179.540 2917.930 181.540 ;
        RECT 0.065 164.540 2917.930 179.540 ;
        RECT 0.065 162.540 2917.200 164.540 ;
        RECT 0.065 161.140 2917.930 162.540 ;
        RECT 2.800 159.140 2917.930 161.140 ;
        RECT 0.065 144.140 2917.930 159.140 ;
        RECT 0.065 142.140 2917.200 144.140 ;
        RECT 0.065 140.740 2917.930 142.140 ;
        RECT 2.800 138.740 2917.930 140.740 ;
        RECT 0.065 123.740 2917.930 138.740 ;
        RECT 0.065 121.740 2917.200 123.740 ;
        RECT 0.065 120.340 2917.930 121.740 ;
        RECT 2.800 118.340 2917.930 120.340 ;
        RECT 0.065 103.340 2917.930 118.340 ;
        RECT 0.065 101.340 2917.200 103.340 ;
        RECT 0.065 99.940 2917.930 101.340 ;
        RECT 2.800 97.940 2917.930 99.940 ;
        RECT 0.065 82.940 2917.930 97.940 ;
        RECT 0.065 80.940 2917.200 82.940 ;
        RECT 0.065 79.540 2917.930 80.940 ;
        RECT 2.800 77.540 2917.930 79.540 ;
        RECT 0.065 62.540 2917.930 77.540 ;
        RECT 0.065 60.540 2917.200 62.540 ;
        RECT 0.065 59.140 2917.930 60.540 ;
        RECT 2.800 57.140 2917.930 59.140 ;
        RECT 0.065 42.140 2917.930 57.140 ;
        RECT 0.065 40.140 2917.200 42.140 ;
        RECT 0.065 38.740 2917.930 40.140 ;
        RECT 2.800 36.740 2917.930 38.740 ;
        RECT 0.065 21.740 2917.930 36.740 ;
        RECT 0.065 19.740 2917.200 21.740 ;
        RECT 0.065 18.340 2917.930 19.740 ;
        RECT 2.800 16.340 2917.930 18.340 ;
        RECT 0.065 1.340 2917.930 16.340 ;
        RECT 0.065 0.175 2917.200 1.340 ;
      LAYER met4 ;
        RECT 15.935 16.495 27.170 3499.105 ;
        RECT 31.070 16.495 45.770 3499.105 ;
        RECT 49.670 16.495 64.370 3499.105 ;
        RECT 68.270 16.495 82.970 3499.105 ;
        RECT 86.870 16.495 101.570 3499.105 ;
        RECT 105.470 16.495 120.170 3499.105 ;
        RECT 124.070 16.495 138.770 3499.105 ;
        RECT 142.670 16.495 188.570 3499.105 ;
        RECT 192.470 16.495 207.170 3499.105 ;
        RECT 211.070 16.495 225.770 3499.105 ;
        RECT 229.670 16.495 244.370 3499.105 ;
        RECT 248.270 16.495 262.970 3499.105 ;
        RECT 266.870 16.495 281.570 3499.105 ;
        RECT 285.470 16.495 300.170 3499.105 ;
        RECT 304.070 16.495 318.770 3499.105 ;
        RECT 322.670 16.495 368.570 3499.105 ;
        RECT 372.470 16.495 387.170 3499.105 ;
        RECT 391.070 16.495 405.770 3499.105 ;
        RECT 409.670 16.495 424.370 3499.105 ;
        RECT 428.270 16.495 442.970 3499.105 ;
        RECT 446.870 16.495 461.570 3499.105 ;
        RECT 465.470 16.495 480.170 3499.105 ;
        RECT 484.070 16.495 498.770 3499.105 ;
        RECT 502.670 16.495 548.570 3499.105 ;
        RECT 552.470 16.495 567.170 3499.105 ;
        RECT 571.070 16.495 585.770 3499.105 ;
        RECT 589.670 16.495 604.370 3499.105 ;
        RECT 608.270 16.495 622.970 3499.105 ;
        RECT 626.870 16.495 641.570 3499.105 ;
        RECT 645.470 16.495 660.170 3499.105 ;
        RECT 664.070 16.495 678.770 3499.105 ;
        RECT 682.670 16.495 728.570 3499.105 ;
        RECT 732.470 16.495 747.170 3499.105 ;
        RECT 751.070 16.495 765.770 3499.105 ;
        RECT 769.670 16.495 784.370 3499.105 ;
        RECT 788.270 16.495 802.970 3499.105 ;
        RECT 806.870 16.495 821.570 3499.105 ;
        RECT 825.470 16.495 840.170 3499.105 ;
        RECT 844.070 16.495 858.770 3499.105 ;
        RECT 862.670 16.495 908.570 3499.105 ;
        RECT 912.470 16.495 927.170 3499.105 ;
        RECT 931.070 16.495 945.770 3499.105 ;
        RECT 949.670 16.495 964.370 3499.105 ;
        RECT 968.270 16.495 982.970 3499.105 ;
        RECT 986.870 16.495 1001.570 3499.105 ;
        RECT 1005.470 16.495 1020.170 3499.105 ;
        RECT 1024.070 16.495 1038.770 3499.105 ;
        RECT 1042.670 16.495 1088.570 3499.105 ;
        RECT 1092.470 16.495 1107.170 3499.105 ;
        RECT 1111.070 16.495 1125.770 3499.105 ;
        RECT 1129.670 16.495 1144.370 3499.105 ;
        RECT 1148.270 16.495 1162.970 3499.105 ;
        RECT 1166.870 16.495 1181.570 3499.105 ;
        RECT 1185.470 16.495 1200.170 3499.105 ;
        RECT 1204.070 16.495 1218.770 3499.105 ;
        RECT 1222.670 16.495 1268.570 3499.105 ;
        RECT 1272.470 16.495 1287.170 3499.105 ;
        RECT 1291.070 16.495 1305.770 3499.105 ;
        RECT 1309.670 16.495 1324.370 3499.105 ;
        RECT 1328.270 16.495 1342.970 3499.105 ;
        RECT 1346.870 16.495 1361.570 3499.105 ;
        RECT 1365.470 16.495 1380.170 3499.105 ;
        RECT 1384.070 16.495 1398.770 3499.105 ;
        RECT 1402.670 16.495 1448.570 3499.105 ;
        RECT 1452.470 16.495 1467.170 3499.105 ;
        RECT 1471.070 16.495 1485.770 3499.105 ;
        RECT 1489.670 16.495 1504.370 3499.105 ;
        RECT 1508.270 16.495 1522.970 3499.105 ;
        RECT 1526.870 16.495 1541.570 3499.105 ;
        RECT 1545.470 16.495 1560.170 3499.105 ;
        RECT 1564.070 16.495 1578.770 3499.105 ;
        RECT 1582.670 16.495 1628.570 3499.105 ;
        RECT 1632.470 16.495 1647.170 3499.105 ;
        RECT 1651.070 16.495 1665.770 3499.105 ;
        RECT 1669.670 16.495 1684.370 3499.105 ;
        RECT 1688.270 16.495 1702.970 3499.105 ;
        RECT 1706.870 16.495 1721.570 3499.105 ;
        RECT 1725.470 16.495 1740.170 3499.105 ;
        RECT 1744.070 16.495 1758.770 3499.105 ;
        RECT 1762.670 16.495 1808.570 3499.105 ;
        RECT 1812.470 16.495 1827.170 3499.105 ;
        RECT 1831.070 16.495 1845.770 3499.105 ;
        RECT 1849.670 16.495 1864.370 3499.105 ;
        RECT 1868.270 16.495 1882.970 3499.105 ;
        RECT 1886.870 16.495 1901.570 3499.105 ;
        RECT 1905.470 16.495 1920.170 3499.105 ;
        RECT 1924.070 16.495 1938.770 3499.105 ;
        RECT 1942.670 16.495 1988.570 3499.105 ;
        RECT 1992.470 16.495 2007.170 3499.105 ;
        RECT 2011.070 16.495 2025.770 3499.105 ;
        RECT 2029.670 16.495 2044.370 3499.105 ;
        RECT 2048.270 16.495 2062.970 3499.105 ;
        RECT 2066.870 16.495 2081.570 3499.105 ;
        RECT 2085.470 16.495 2100.170 3499.105 ;
        RECT 2104.070 16.495 2118.770 3499.105 ;
        RECT 2122.670 16.495 2168.570 3499.105 ;
        RECT 2172.470 16.495 2187.170 3499.105 ;
        RECT 2191.070 16.495 2205.770 3499.105 ;
        RECT 2209.670 16.495 2224.370 3499.105 ;
        RECT 2228.270 16.495 2242.970 3499.105 ;
        RECT 2246.870 16.495 2261.570 3499.105 ;
        RECT 2265.470 16.495 2280.170 3499.105 ;
        RECT 2284.070 16.495 2298.770 3499.105 ;
        RECT 2302.670 16.495 2348.570 3499.105 ;
        RECT 2352.470 16.495 2367.170 3499.105 ;
        RECT 2371.070 16.495 2385.770 3499.105 ;
        RECT 2389.670 16.495 2404.370 3499.105 ;
        RECT 2408.270 16.495 2422.970 3499.105 ;
        RECT 2426.870 16.495 2441.570 3499.105 ;
        RECT 2445.470 16.495 2460.170 3499.105 ;
        RECT 2464.070 16.495 2478.770 3499.105 ;
        RECT 2482.670 16.495 2528.570 3499.105 ;
        RECT 2532.470 16.495 2547.170 3499.105 ;
        RECT 2551.070 16.495 2565.770 3499.105 ;
        RECT 2569.670 16.495 2584.370 3499.105 ;
        RECT 2588.270 16.495 2602.970 3499.105 ;
        RECT 2606.870 16.495 2621.570 3499.105 ;
        RECT 2625.470 16.495 2640.170 3499.105 ;
        RECT 2644.070 16.495 2658.770 3499.105 ;
        RECT 2662.670 16.495 2708.570 3499.105 ;
        RECT 2712.470 16.495 2727.170 3499.105 ;
        RECT 2731.070 16.495 2745.770 3499.105 ;
        RECT 2749.670 16.495 2764.370 3499.105 ;
        RECT 2768.270 16.495 2782.970 3499.105 ;
        RECT 2786.870 16.495 2801.570 3499.105 ;
        RECT 2805.470 16.495 2820.170 3499.105 ;
        RECT 2824.070 16.495 2838.770 3499.105 ;
        RECT 2842.670 16.495 2888.570 3499.105 ;
        RECT 2892.470 16.495 2905.985 3499.105 ;
  END
END user_analog_project_wrapper
END LIBRARY

